// de1_soc_hex_display.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module de1_soc_hex_display (
		input  wire        hex_0_clk_clk,                    //                 hex_0_clk.clk
		output wire [6:0]  hex_0_external_connection_export, // hex_0_external_connection.export
		input  wire        hex_0_reset_reset_n,              //               hex_0_reset.reset_n
		input  wire [1:0]  hex_0_s1_address,                 //                  hex_0_s1.address
		input  wire        hex_0_s1_write_n,                 //                          .write_n
		input  wire [31:0] hex_0_s1_writedata,               //                          .writedata
		input  wire        hex_0_s1_chipselect,              //                          .chipselect
		output wire [31:0] hex_0_s1_readdata,                //                          .readdata
		input  wire        hex_1_clk_clk,                    //                 hex_1_clk.clk
		output wire [6:0]  hex_1_external_connection_export, // hex_1_external_connection.export
		input  wire        hex_1_reset_reset_n,              //               hex_1_reset.reset_n
		input  wire [1:0]  hex_1_s1_address,                 //                  hex_1_s1.address
		input  wire        hex_1_s1_write_n,                 //                          .write_n
		input  wire [31:0] hex_1_s1_writedata,               //                          .writedata
		input  wire        hex_1_s1_chipselect,              //                          .chipselect
		output wire [31:0] hex_1_s1_readdata,                //                          .readdata
		input  wire        hex_2_clk_clk,                    //                 hex_2_clk.clk
		output wire [6:0]  hex_2_external_connection_export, // hex_2_external_connection.export
		input  wire        hex_2_reset_reset_n,              //               hex_2_reset.reset_n
		input  wire [1:0]  hex_2_s1_address,                 //                  hex_2_s1.address
		input  wire        hex_2_s1_write_n,                 //                          .write_n
		input  wire [31:0] hex_2_s1_writedata,               //                          .writedata
		input  wire        hex_2_s1_chipselect,              //                          .chipselect
		output wire [31:0] hex_2_s1_readdata,                //                          .readdata
		input  wire        hex_3_clk_clk,                    //                 hex_3_clk.clk
		output wire [6:0]  hex_3_external_connection_export, // hex_3_external_connection.export
		input  wire        hex_3_reset_reset_n,              //               hex_3_reset.reset_n
		input  wire [1:0]  hex_3_s1_address,                 //                  hex_3_s1.address
		input  wire        hex_3_s1_write_n,                 //                          .write_n
		input  wire [31:0] hex_3_s1_writedata,               //                          .writedata
		input  wire        hex_3_s1_chipselect,              //                          .chipselect
		output wire [31:0] hex_3_s1_readdata,                //                          .readdata
		input  wire        hex_4_clk_clk,                    //                 hex_4_clk.clk
		output wire [6:0]  hex_4_external_connection_export, // hex_4_external_connection.export
		input  wire        hex_4_reset_reset_n,              //               hex_4_reset.reset_n
		input  wire [1:0]  hex_4_s1_address,                 //                  hex_4_s1.address
		input  wire        hex_4_s1_write_n,                 //                          .write_n
		input  wire [31:0] hex_4_s1_writedata,               //                          .writedata
		input  wire        hex_4_s1_chipselect,              //                          .chipselect
		output wire [31:0] hex_4_s1_readdata,                //                          .readdata
		input  wire        hex_5_clk_clk,                    //                 hex_5_clk.clk
		output wire [6:0]  hex_5_external_connection_export, // hex_5_external_connection.export
		input  wire        hex_5_reset_reset_n,              //               hex_5_reset.reset_n
		input  wire [1:0]  hex_5_s1_address,                 //                  hex_5_s1.address
		input  wire        hex_5_s1_write_n,                 //                          .write_n
		input  wire [31:0] hex_5_s1_writedata,               //                          .writedata
		input  wire        hex_5_s1_chipselect,              //                          .chipselect
		output wire [31:0] hex_5_s1_readdata                 //                          .readdata
	);

	de1_soc_hex_display_hex_0 hex_0 (
		.clk        (hex_0_clk_clk),                    //                 clk.clk
		.reset_n    (hex_0_reset_reset_n),              //               reset.reset_n
		.address    (hex_0_s1_address),                 //                  s1.address
		.write_n    (hex_0_s1_write_n),                 //                    .write_n
		.writedata  (hex_0_s1_writedata),               //                    .writedata
		.chipselect (hex_0_s1_chipselect),              //                    .chipselect
		.readdata   (hex_0_s1_readdata),                //                    .readdata
		.out_port   (hex_0_external_connection_export)  // external_connection.export
	);

	de1_soc_hex_display_hex_0 hex_1 (
		.clk        (hex_1_clk_clk),                    //                 clk.clk
		.reset_n    (hex_1_reset_reset_n),              //               reset.reset_n
		.address    (hex_1_s1_address),                 //                  s1.address
		.write_n    (hex_1_s1_write_n),                 //                    .write_n
		.writedata  (hex_1_s1_writedata),               //                    .writedata
		.chipselect (hex_1_s1_chipselect),              //                    .chipselect
		.readdata   (hex_1_s1_readdata),                //                    .readdata
		.out_port   (hex_1_external_connection_export)  // external_connection.export
	);

	de1_soc_hex_display_hex_0 hex_2 (
		.clk        (hex_2_clk_clk),                    //                 clk.clk
		.reset_n    (hex_2_reset_reset_n),              //               reset.reset_n
		.address    (hex_2_s1_address),                 //                  s1.address
		.write_n    (hex_2_s1_write_n),                 //                    .write_n
		.writedata  (hex_2_s1_writedata),               //                    .writedata
		.chipselect (hex_2_s1_chipselect),              //                    .chipselect
		.readdata   (hex_2_s1_readdata),                //                    .readdata
		.out_port   (hex_2_external_connection_export)  // external_connection.export
	);

	de1_soc_hex_display_hex_0 hex_3 (
		.clk        (hex_3_clk_clk),                    //                 clk.clk
		.reset_n    (hex_3_reset_reset_n),              //               reset.reset_n
		.address    (hex_3_s1_address),                 //                  s1.address
		.write_n    (hex_3_s1_write_n),                 //                    .write_n
		.writedata  (hex_3_s1_writedata),               //                    .writedata
		.chipselect (hex_3_s1_chipselect),              //                    .chipselect
		.readdata   (hex_3_s1_readdata),                //                    .readdata
		.out_port   (hex_3_external_connection_export)  // external_connection.export
	);

	de1_soc_hex_display_hex_0 hex_4 (
		.clk        (hex_4_clk_clk),                    //                 clk.clk
		.reset_n    (hex_4_reset_reset_n),              //               reset.reset_n
		.address    (hex_4_s1_address),                 //                  s1.address
		.write_n    (hex_4_s1_write_n),                 //                    .write_n
		.writedata  (hex_4_s1_writedata),               //                    .writedata
		.chipselect (hex_4_s1_chipselect),              //                    .chipselect
		.readdata   (hex_4_s1_readdata),                //                    .readdata
		.out_port   (hex_4_external_connection_export)  // external_connection.export
	);

	de1_soc_hex_display_hex_0 hex_5 (
		.clk        (hex_5_clk_clk),                    //                 clk.clk
		.reset_n    (hex_5_reset_reset_n),              //               reset.reset_n
		.address    (hex_5_s1_address),                 //                  s1.address
		.write_n    (hex_5_s1_write_n),                 //                    .write_n
		.writedata  (hex_5_s1_writedata),               //                    .writedata
		.chipselect (hex_5_s1_chipselect),              //                    .chipselect
		.readdata   (hex_5_s1_readdata),                //                    .readdata
		.out_port   (hex_5_external_connection_export)  // external_connection.export
	);

endmodule
