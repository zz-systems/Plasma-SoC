---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"8E3CAF273C14AC2C008C3C00088C3C24088C3C3C000000000003273C0003273C",
INIT_01 => X"3CAF3C2727038F8F8F240824AC3C3CAE1000162A0C24AC24AFAE3C00243CAF24",
INIT_02 => X"1002008E00162402122400300C008C3C001402263CAF14AFAFAFAF00243C8E8C",
INIT_03 => X"3C8E3CAF27001030008C3C27038F8F8F8F8F8FA0AE241200008EA01024AC243C",
INIT_04 => X"27083C8F8F000C8E240C3C8E240C008E240C3C8E240C008E000C8C8E3C240CAF",
INIT_05 => X"AF8CAF3C2727038FA28F8FA200932410A20012932A0CAF020027AF00AF270003",
INIT_06 => X"8F8E8F8F8F8F00021424240C000002168EAC0C0000AF24AF268E3CAF00021624",
INIT_07 => X"AC8C243C243C243C241400AC243C243C241400AC243C243C273C273C00270800",
INIT_08 => X"AFAFAFAFAFAFAFAFAFAF2308000C000C24142400AC8C243C243C243C24142400",
INIT_09 => X"8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F000CAF00AF00AF2340AFAFAFAFAFAFAFAF",
INIT_0A => X"248C0003001030008C0003001030008C0040034040033423038F038F8F8F8F8F",
INIT_0B => X"ACAC3C0010240CAFAF00AF270003AC00248C0003AC34008C0003AC00008CAC34",
INIT_0C => X"3C14020C2424103C3C14020C24AE1024AE243C3C14020C2424103C3C14020C24",
INIT_0D => X"2410AE243C3C14020C242410AE243C3C14020C242410AE3C3C14020C2424103C",
INIT_0E => X"AF3CAF2700000010000CAF2700000027038F8F028F00020C2410AE3C14020C24",
INIT_0F => X"16263C0C0202000010008E00120014020210028E24243C000026AFAFAFAFAFAF",
INIT_10 => X"003C0C3002003C0C02AC0024AFAF00240030AF3C2727038F8F8F8F8F8F8F8F26",
INIT_11 => X"10248C3C0024240010AC03ACACAC24AC3C00343C0024243C27083C308F028F8F",
INIT_12 => X"ACACACAC008C8C000300108CAC10ACACAC008CACAC240024142C001400008C00",
INIT_13 => X"1000108C008CACACACAC8C00108CAC10ACACAC8C001100001024248C3C100003",
INIT_14 => X"001000000000000300108C000000ACACACAC008C8CAC2400008C001400008C24",
INIT_15 => X"308CAC0000008C240003AC00008CAC0000248C000300248C00000000032410AC",
INIT_16 => X"000003AC0000308CAC0000008C240003AC0000308CAC0000008C240003AC0000",
INIT_17 => X"0003AC00341024108C0003AC0000308CAC00248C0003AC340003ACAC340003AC",
INIT_18 => X"0003AC00008CAC34248C0003AC00248C0003AC34008C000800080008000003AC",
INIT_19 => X"1624ACACACAC0010000C2400AF12AFAFAF8CAF2700000003AC00008CAC34248C",
INIT_1A => X"0CAE14240C00100010322424001024AE24AEAE243C16240010AEAE24AEAE243C",
INIT_1B => X"000CAFAFAF2727038F8F8F8F028FAEAE24AE10240C0012001232AEAE24001002",
INIT_1C => X"8F8F27088F028F8F2400102410020C243C10020C243C2410020C243C10008C00",
INIT_1D => X"10008100AF000027000300AC242403A0AC24001000008C8C3010008C2703008F",
INIT_1E => X"24000390AC24001000008C8C0010008C2703008F0000100010008D00250C0130",
INIT_1F => X"8C0010008CAC00008C0010008C241400100014008CAC0010008C2414000300AC",
INIT_20 => X"14AFAFAF248C278C0003AC0000008C0010008CAC0000008C0010008C00140010",
INIT_21 => X"10248C008E000CAFAF270010260C8C928E001002008E8C270800008F028F8F00",
INIT_22 => X"000024000CAF270003241000100080000027088F028F000C8E000C8E000C8E00",
INIT_23 => X"10A110002400002400001524000000002703008FA01024A02480800010000000",
INIT_24 => X"248024000000033403000030302410241000140080800008A000A12424000400",
INIT_25 => X"8FAE8F000C00AFAFAF2727038F8E8F000CAFAF2700000008000800080003A014",
INIT_26 => X"AFAFAF272703308F8F8E000CAFAF2727038F8F00AE8F000C30AFAFAF2727038F",
INIT_27 => X"0027038F8F8F8F8F8F0010AE020C9226AE020C00140010008224240000AFAFAF",
INIT_28 => X"3C3C240C240C243C240C243C240C243C240C243C240C243CAF0CAFAF2400273C",
INIT_29 => X"0C36240C36240C263C3C0C3C0C3C0CAC0C3C3C240C243C3CAE0C263C240C243C",
INIT_2A => X"360C360C24240C36240C26240C36240C36340C263C240C36240C36240C263C24",
INIT_2B => X"544F4C494F4C4921544953412703008F8F8F240C243C3C240C3C8C3C240C3C8E",
INIT_2C => X"7463640074636400746364007463640030300D4D6C0D006C646477307564723A",
INIT_2D => X"0003273C0003273C000000000000000000000000000000007230676400696400",
INIT_2E => X"0000006569616743002E6161742E612E65455443646C2E2E6E61730000000F41",
INIT_2F => X"646C2E2E6E61730000000F410003273C0003273C000000000000000000000000",
INIT_30 => X"0000000000000000000000000000006569616743002E6161742E612E65455443",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"2311B1BD0440644400620300004402A5004405020000000000405A1A00405A1A",
INIT_01 => X"12B202BDBDE0B0B1BF8400A54005022000000010008443A5BF3002627005B002",
INIT_02 => X"4003008300620240620213A5000544024060233111B080B1B3B4BF6242024345",
INIT_03 => X"050410B0BD004042004202BDE0B0B1B2B3B4BF53434320510042620002446402",
INIT_04 => X"BD0004B0BF000004A500050405000004A5000504050000040000450402A500BF",
INIT_05 => X"B150B002BDBDE0B002B1BF0300A30200020020A23100BF2080A5B0A0B1BD00E0",
INIT_06 => X"B244B0B1B3BF0705A0058400000771204443000000BF84B3034412B207112011",
INIT_07 => X"A3C38404A505C606A560A4A08404A505A560A4A08404A505BD1D9C1C00BD0000",
INIT_08 => X"AAA9A8A7A6A5A4A3A2A1BD0000000000A560C6A4A3C38404A505C606A560C6A4",
INIT_09 => X"AFAEADACABAAA9A8A7A6A5A4A3A2A10000BB00BB00BA5A1ABFB9B8AFAEADACAB",
INIT_0A => X"038200E0004042008200E000404200820084E0029B401BBD60BB60BBBABFB9B8",
INIT_0B => X"40400540400400BFB080B1BD00E08243038200E08242008200E0824300828242",
INIT_0C => X"05402000A542000205402000A502000202420205402000A542000205402000A5",
INIT_0D => X"020002420205402000A5020002420205402000A50200020205402000A5420002",
INIT_0E => X"B611B1BD000000000000BFBD000000BDE0B0B100BF00000002000202402000A5",
INIT_0F => X"14100400007240004000220040004053424016A2141615000031B2BFB0B3B4B5",
INIT_10 => X"100400C6201004002044A006B0BF624211B1B102BDBDE0B0B1B2B3B4B5B6BF31",
INIT_11 => X"62424302828402008082E043436283430462630343420302BD0004C6B120B0BF",
INIT_12 => X"606085A400656400E00000636600C3C486006464C5A54462C0A6A4C0A4006500",
INIT_13 => X"600045460062468287E6E2000042E600878246470000C2E047678662038000E0",
INIT_14 => X"00668680800600E00000C6C04060404087E400444764848700470047E4006467",
INIT_15 => X"C682824302A2830200E085A2058283A3A20283A2E0A3038200000000E0630065",
INIT_16 => X"0000E085A2A6C682824302A2830200E085A2A6C682824302A2830200E085A2A6",
INIT_17 => X"00E08243420003A08200E085A205A5828243038200E085A500E08582A200E085",
INIT_18 => X"00E0824300828242038200E08243038200E0824200820000000000000000E085",
INIT_19 => X"6202404040524040A0000480B060B1B2BF93B3BD000000E08243008282420382",
INIT_1A => X"0002400400004000602302120000120202020242026202000000020202024202",
INIT_1B => X"A000BFB0B1BDBDE0B0B1B2B300BF020303024004000040002031020303000000",
INIT_1C => X"B1BFBD00B120B0BF05000005400000A505400000A50505400000A50540004240",
INIT_1D => X"A0000500BFA080BD00E000820202E0C582C20060C2438683A5400082BDE000B0",
INIT_1E => X"0200E0A282A20060A243858300400082BDE000BF000000E0400022E2080020A5",
INIT_1F => X"8200400082824500820040008202C2000000400082824540008202C000E00082",
INIT_20 => X"62B1BFB00243BD8200E08545A30083004000828243A300830040008200C24500",
INIT_21 => X"62024300028000BFB0BD00003100442502004022000291BD000000B000B1BF80",
INIT_22 => X"8082428000BFBD44E04200006000438000BD00B000BF00000400000400000400",
INIT_23 => X"00074000E700A3C30749200900436404BDE000BF440042666346640080864565",
INIT_24 => X"63A4A5808000E042E002434263A5008440004300A382A00060A302C302A38160",
INIT_25 => X"B111BF8000A0B0B1BFBDBDE0B002BF8000B0BFBD000000000000000000E06480",
INIT_26 => X"B1B2B3BDBDE042B0BF028000BFB0BDBDE0B0B10011BF8000B1B0B1BFBDBDE0B0",
INIT_27 => X"00BDE0B0B1B2B3B4BF000034200014103320000052004000021312A080B4BFB0",
INIT_28 => X"040504008400050484000504840005048400050484000504B000B1BF8400BD04",
INIT_29 => X"0004050004A5000405040004000400620004038400A50405220004118400A510",
INIT_2A => X"0400040005050004050004050004050004A5000405050004050004A500040505",
INIT_2B => X"694645524E45520D494F5343BDE000B0B1BF8400A50405A500054402A5000524",
INIT_2C => X"656F6500656F6500656F6500656F65003A300A416C0A00616965000061657720",
INIT_2D => X"00405A1A00405A1A000000000000000000000000000000000000706500726500",
INIT_2E => X"0000007362746E4B536274006469747278004154006462676F62742E07016700",
INIT_2F => X"006462676F62742E0701670000405A1A00405A1A000000000000000000000000",
INIT_30 => X"0000000000000000000000000000007362746E4B536274006469747278004154",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"170000FF00001700001700000417001503170000000000000000040000000300",
INIT_01 => X"000020FF00000000001704150400201700000000041704150017201800000000",
INIT_02 => X"00100016000000A000009E00039E170080001817000000000000002016001601",
INIT_03 => X"00170000FF000000000040000000000000000000160000880016FF000016FF00",
INIT_04 => X"0003400000000417160300170003301717030017000330170003161700150300",
INIT_05 => X"00170000FF000000000000000000000000000000000400208000008800FF0000",
INIT_06 => X"0016000000000000000E00002800000016170098280000000016000000000000",
INIT_07 => X"000016001600160000FF18001600160000FF1800170016001900160000000028",
INIT_08 => X"00000000000000000000FF010001000200FF0018000016001600160000FF0018",
INIT_09 => X"000000000000000000000000000000000100D800D800FF700000000000000000",
INIT_0A => X"FF00000000FF000000000000FF00000000600060600000000000000000000000",
INIT_0B => X"0000008000000200008800FF00000010FF000000000000000000001000000000",
INIT_0C => X"000020041603FF20000020041600000000032000002004160300200000200416",
INIT_0D => X"00FF000120000020041600FF000420000020041600FF0020000020041603FF20",
INIT_0E => X"000000FF000000FF000500FF00000000000000100080200200FF004000200416",
INIT_0F => X"FF0020022898F800000000000000001090009000000020988017000000000000",
INIT_10 => X"3420020028342002280080000000101718000000FF0000000000000000000000",
INIT_11 => X"001616002000FF1000160000000016000018FF001019FF000002200000280000",
INIT_12 => X"00000000000000100000FF00000000000000000000FF30000000280030000000",
INIT_13 => X"00000000181600FFFF000000FF000000FFFF0000000040280016FF1600000000",
INIT_14 => X"000030181030000000FF00101810000000000000000000200000000038000000",
INIT_15 => X"000000101010000000000028280000182800001000280000000000000000FF00",
INIT_16 => X"0000000028280000001010100000000000282800000010101000000000002828",
INIT_17 => X"000000100000FF0000000000282800000010FF00000000000000000000000000",
INIT_18 => X"0000001000000000FF0000000010FF0000000000000000010001000100000000",
INIT_19 => X"00000000000080008804009000000000000000FF00000000001000000000FF00",
INIT_1A => X"0400000004000000000000001000000000000001200000900000000000000040",
INIT_1B => X"8001000000FF000000000000100000000000FF00040000000000000000800020",
INIT_1C => X"0000000300200000000000000020041600002004160000002004160000000088",
INIT_1D => X"00000038004048FF000010000000000000001000181000000000000000001000",
INIT_1E => X"000000000000100018100000000000000000000010000010FF00003800032000",
INIT_1F => X"0000000000001000000000000000000000000000000010000000000000001000",
INIT_20 => X"000000000000FF00000000282800000000000000101800000000000000002800",
INIT_21 => X"000000000080040000FF00FF000400000000FF10000000000328300020000080",
INIT_22 => X"1810FF280400FF100000FF000000001000000400200000040000040000040000",
INIT_23 => X"FFFF001000384000000000003010101F0000000000FFFFFF0000000000203020",
INIT_24 => X"00FF001810100000001010000000FF0000000000000020040018000000180030",
INIT_25 => X"000000800188000000FF000000000080010000FF00000002000200020000FFFF",
INIT_26 => X"000000FF00000000000080010000FF00000000100000800100000000FF000000",
INIT_27 => X"00000000000000000000FF002001FF0000200100000000000000008088000000",
INIT_28 => X"000000010002000000020000000200000102000002020000000200000028FF00",
INIT_29 => X"0203000203120203004001400340031701400016031600001701010016031620",
INIT_2A => X"0201020300000202000202000203000203A10203000002030002035E02030000",
INIT_2B => X"6D4644432044430A4F4C20430000100000001604160000160400160016030017",
INIT_2C => X"72757600727576007275760072757600303A00496F4800797376000072760000",
INIT_2D => X"0000040000000300000016160000161600001616000016160000697600637600",
INIT_2E => X"00000000757475005473612E616E616F742E424F562D756E7400727304006E00",
INIT_2F => X"562D756E7400727304006E000000040000000300000000000000000000000000",
INIT_30 => X"00000000000000000000000000000000757475005473612E616E616F742E424F",
INIT_31 => X"0000161500000000000000150000000000000000000017000000000000000000",
INIT_32 => X"0000000017160000000000000000171600000000000000001716000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000002171700000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"200018E000161C01001C0000181400D0B8140000000000000008540000089000",
INIT_01 => X"001800D8200814181C009BF008000020070009089B0008E41C20000401001401",
INIT_02 => X"0D2B00C0000B7F25040803FFA4001400251E2B00001023141C20242BE000C008",
INIT_03 => X"00100010E800260100040028081014181C202400C001032B00C0FF0820C0FF00",
INIT_04 => X"1816001014001810E0B8001020E4251000B8001010E4251000B8C41000FCB814",
INIT_05 => X"18181400D828081C0020240100113004010004100A70242525101C2520D80008",
INIT_06 => X"1CC4141820240D1A021003A2100D1A02C418A2121024062001C4001C0D1A023C",
INIT_07 => X"0000E000C000A00004FD2A00E000E00004FD2A00B000E000B000E0000028A212",
INIT_08 => X"34302C2824201C181410981400D4002804FB042A0000E000E000C00004FB042A",
INIT_09 => X"4844403C3834302C2824201C18141000DC60125C1058FC0054504C4844403C38",
INIT_0A => X"FE00000800FC020004000800FC01000400000800000801681360115C5854504C",
INIT_0B => X"040000254F08371C142518E000080024FD000008000200000008002400000001",
INIT_0C => X"0004258A7420F5000004258A640439010010000007258A540008000004258A44",
INIT_0D => X"05D20000000006258A0804DC0000000006258A9003E600000005258A8430ED00",
INIT_0E => X"280014D0000000FF000014E800000020081418251C25256207CA000004258A18",
INIT_0F => X"EC0100AD25250900060000000A000C2424120408200100252530182C101C2024",
INIT_10 => X"4200C501250200B825002501141C2130801F1800E030081014181C2024282C04",
INIT_11 => X"17D0D0002403FC2528D008040004D0080023F47F24B3FC0020D200011825141C",
INIT_12 => X"00040004000004250800E900000604000400000808F4210C1104230F2B000800",
INIT_13 => X"13001A0025D000F8F4040400F3000009F8F4040400072B250DD0F4D000350008",
INIT_14 => X"000421252580000800E600252525000400040004000810210008000E2100080C",
INIT_15 => X"011818242704180100081024271010250401102408040100000000000804FC00",
INIT_16 => X"0000081C2504011C1C2427041C01000814250401141424270414010008182504",
INIT_17 => X"000800240402FB030000080025C007000024C70000080002000800000100080C",
INIT_18 => X"0008002400000010EF0000080024F700000800080000006E0068005E0000080C",
INIT_19 => X"09071C080400252825A42025142E181C240420D800000008002400000020DF00",
INIT_1A => X"A6040540A4000C000E01010125030114010C0408000905250A14184010080800",
INIT_1B => X"25741C1418E0280814181C20252410184008F140A40008000A020C1440251025",
INIT_1C => X"181C202C1825141C0200080104258A9C0008258A1400030F258A04001A000425",
INIT_1D => X"0B000025142525E80008251C02010800100125092B211018FF0C000820082514",
INIT_1E => X"020008000C0125042B210C14000C00041808001425000225F5001C2101A425FF",
INIT_1F => X"0C00180004102100100005000802100026002600041021020008010C0008251C",
INIT_20 => X"09181C140704E00000080C212100140006000410212100180006000800132114",
INIT_21 => X"070704000025181410E800F501C300000000F32B00100820E425251425181C25",
INIT_22 => X"2521FF255014E8230801FB00030000250018A610251400A60000A60800A60400",
INIT_23 => X"F5FF0312301021010D1A020A252326C31808001401F5FFFF01000000082A2323",
INIT_24 => X"01FF01252525080108232BFFFF01F8010900050000002559002100022D210525",
INIT_25 => X"18081C25502514181CE0180810081425571014E80000009A006200370008FFFC",
INIT_26 => X"14181CD81808FF10140825571410E82008141825081C2550FF14181CE0200814",
INIT_27 => X"0028081014181C202400F1082550FF010825500004000D00000D0A2525202410",
INIT_28 => X"0000014C300B1F00440B0800540B0700D40B0600EC0B0200140B181CF025E000",
INIT_29 => X"E80008E300D0E0001300500020000A10680000187A14000014680000087A0400",
INIT_2A => X"006800000101F70004EC000CE82008E32020E020070CE81008E31010E0105F0C",
INIT_2B => X"65002020002020004E41564520082514181CE09B400000389B00C40028B80014",
INIT_2C => X"336E2F00326E2F00316E2F00306E2F003030004E20650030702F0000742F0000",
INIT_2D => X"00085400000890000000D0D0000038E00000D0D0000038E000006F2F00302F00",
INIT_2E => X"0000000074722E2E417300647469006400744C5245696975652E746801007500",
INIT_2F => X"45696975652E7468010075000008540000089000A00002070B00000000000000",
INIT_30 => X"A00002070B000000000000000000000074722E2E417300647469006400744C52",
INIT_31 => X"00D070D032013000100000A0D03007012A0001000020600000011E0004000024",
INIT_32 => X"100000D060E0030848001000002040C0030142000100002040A0030838010400",
INIT_33 => X"000000000000000000000000000000000000000053000100000060B003084D00",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic