---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"8E3CAF273C14AC2C008C3C00088C3C24088C3C3C000000000003273C0003273C",
INIT_01 => X"008C3C27038F8F2408AC8C3C3CAE10001428008E000CAC24AF3C8C0024AE243C",
INIT_02 => X"003C2400340003000327083C8F8F000C8E240C3C8E3C0C3CAF0CAF3C27001030",
INIT_03 => X"241400AC243C243C241400AC243C243C273C273C0000030014008C3CAC24ACAC",
INIT_04 => X"AFAF2308000C000C24142400AC8C243C243C243C24142400AC8C243C243C243C",
INIT_05 => X"200010002000108C3CAF00AF00AF2340AFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAF",
INIT_06 => X"8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F0008ACAC3C00208F230CAF0008",
INIT_07 => X"008CAC34248C0003001030008C0003001030008C0040034040033423038F038F",
INIT_08 => X"0003AC3C3400033C13008C00243C00240003AC00248C0003AC34008C0003AC00",
INIT_09 => X"03AC00308CAC00008CAC0030008CAC00008CAC00008C3CAC00243C0024002430",
INIT_0A => X"00008C0010248C3C0024240010AC03ACACAC24AC3C00343C0024243C00000000",
INIT_0B => X"3C100003ACACACAC008C8C000300108CAC10ACACAC008CACAC240024142C0014",
INIT_0C => X"00008C241000108C008CACACACAC8C00108CAC10ACACAC8C001100001024248C",
INIT_0D => X"0003ACAC340003AC0000000300108C000000ACACACAC008C8CAC2400008C0014",
INIT_0E => X"0003AC00008CAC34248C0003AC00248C0003AC34008C0008000800080003AC34",
INIT_0F => X"1624ACACACAC0010000C2400AF12AFAFAF8CAF2700000003AC00008CAC34248C",
INIT_10 => X"27038F8F8F8F028FAE0010020CAE14240C001232AEAE10240C001032AE10243C",
INIT_11 => X"8F8F2400102410020C243C10020C243C2410020C243C10008C00000CAFAFAF27",
INIT_12 => X"000027000300AC242403A0AC24001000248C3010008C2703008F8F8F27088F02",
INIT_13 => X"8C24140003AC240014008C2703008F0000100010008D00250C013010008100AF",
INIT_14 => X"278C0003AC00008C0010008CAC00008C0010008C001400100014008CAC001000",
INIT_15 => X"0CAFAF270010260C8C928E001002008E8C270800008F028F8F0014AFAFAF248C",
INIT_16 => X"032410001000800000000027088F028F000C8E000C8E000C8E0010248C008E00",
INIT_17 => X"00001524000000002703008FA01024A02480800010000000000024000CAF2700",
INIT_18 => X"03000030302410241000140080800008A000A1242400040010A1100024000024",
INIT_19 => X"2727038F8FAE8F000C00AFAFAF2727038F8E8F000CAFAF270008000800000334",
INIT_1A => X"0000AFAFAFAFAFAF2727038F8E8F000CAFAF2727038F8F00AE8F000C00AFAFAF",
INIT_1B => X"AF00AF27000027038F8F8F8F8F8F0010AE020C8226AE020C0014001000822424",
INIT_1C => X"3C3C14020C242410AE243C3C14020C2424103C3C14020C24ACAC3C0010240CAF",
INIT_1D => X"020C242410AE243C3C14020C242410AE3C3C14020C2424103C3C14020C242410",
INIT_1E => X"AF0CAFAF2424273C00000027038F8F028FAE24AE3C14020C242410AE243C3C14",
INIT_1F => X"0C3C3C240C243C3CAE0C263C240C243C3C3C240C240C243C240C243C240C243C",
INIT_20 => X"0C24360C24260C343C360C24360C24260C243C360C24360C24260C243C3C0CAC",
INIT_21 => X"48006C6464773075647221540A4F4C49004F4C4921544953410010240C8E3C36",
INIT_22 => X"000000000000306764006964007463640074636400746364007463647200496F",
INIT_23 => X"742E612E65455443646C2E2E6E61730000000F410003273C0003273C00000000",
INIT_24 => X"00000000000000000000000000000000000000000000006569616743002E6161",
INIT_25 => X"65455443646C2E2E6E61730000000F410003273C0003273C0000000000000000",
INIT_26 => X"000000000000000000000000000000000000006569616743002E6161742E612E",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"0310B0BD0440644400620300004402A5004405020000000000405A1A00405A1A",
INIT_01 => X"004202BDE0B0BFA5004084050200000040420002000043A5BF02846202026205",
INIT_02 => X"000203820200E000E0BD0004B0BF000004A5000504040010B000BF04BD004042",
INIT_03 => X"A560A4A08404A505A560A4A08404A505BD1D9C1C0000E0004000620343034344",
INIT_04 => X"A2A1BD0000000000A560C6A4A3C38404A505C606A560C6A4A3C38404A505C606",
INIT_05 => X"8406A8C5050006C606BB00BB00BA5A1ABFB9B8AFAEADACABAAA9A8A7A6A5A4A3",
INIT_06 => X"BABFB9B8AFAEADACABAAA9A8A7A6A5A4A3A2A10000C0C5068505A4A500A40000",
INIT_07 => X"00828242038200E0004042008200E000404200820084E0029B401BBD60BB60BB",
INIT_08 => X"00E0430263002003200099448404048400E08243038200E08242008200E08243",
INIT_09 => X"E045A3A54343640544448684054644830344446400440244C2420202424303A2",
INIT_0A => X"A400650062424302828402008082E04343628343046263034342030200000000",
INIT_0B => X"038000E0606085A400656400E00000636600C3C486006464C5A54462C0A6A4C0",
INIT_0C => X"E4006467600045460062468287E6E2000042E600878246470000C2E047678662",
INIT_0D => X"00E08582A200E085000000E00000C6C04060404087E400444764848700470047",
INIT_0E => X"00E0824300828242038200E08243038200E08242008200000000000000E085A5",
INIT_0F => X"6202404040524040A0000480B060B1B2BF93B3BD000000E08243008282420382",
INIT_10 => X"BDE0B0B1B2B300BF020000000002400400002031020240040000402202004202",
INIT_11 => X"B0BF05000005400000A505400000A50505400000A50540004240A000BFB0B1BD",
INIT_12 => X"A080BD00E000820202E0C582C20060C24286A5400082BDE000B0B1BFBD00B120",
INIT_13 => X"8202C000E0820200400082BDE000BF000000E0400022E2080020A5A0000500BF",
INIT_14 => X"BD8200E08545008200400082824500820040008200C200000040008282454000",
INIT_15 => X"00BFB0BD00003100442502004022000291BD000000B000B1BF8062B1BFB00243",
INIT_16 => X"E042000060004380000000BD00B000BF00000400000400000400620243000280",
INIT_17 => X"0749200900436404BDE000BF4400426663466400808645658082428000BFBD44",
INIT_18 => X"E002434263A5008440004300A382A00060A302C302A3816000074000E700A3C3",
INIT_19 => X"BDBDE0B0B111BF8000A0B0B1BFBDBDE0B002BF8000B0BFBD000000000000E042",
INIT_1A => X"A080B4BFB0B1B2B3BDBDE0B002BF8000B0BFBDBDE0B0B10011BF8000A0B0B1BF",
INIT_1B => X"B080B1BD0000BDE0B0B1B2B3B4BF000034200014103320000052004000021312",
INIT_1C => X"0205402000A5020002420205402000A542000205402000A540400540400400BF",
INIT_1D => X"2000A5020002420205402000A50200020205402000A542000205402000A54200",
INIT_1E => X"B000B1BF8405BD04000000BDE0B0B100BF02020202402000A502000242020540",
INIT_1F => X"0004038400A50405220004118400A51004050400840005048400050484000504",
INIT_20 => X"00050400050400A5050400050400050400A5050400050400050400A505040062",
INIT_21 => X"65006169650000616577006500464552004E45520D494F53430000A500240504",
INIT_22 => X"00000000000000706500726500656F6500656F6500656F6500656F6500004E20",
INIT_23 => X"6469747278004154006462676F62742E0701670000405A1A00405A1A00000000",
INIT_24 => X"00000000000000000000000000000000000000000000007362746E4B53627400",
INIT_25 => X"78004154006462676F62742E0701670000405A1A00405A1A0000000000000000",
INIT_26 => X"000000000000000000000000000000000000007362746E4B5362740064697472",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"110000FF00001100001100000211001002110000000000000000020000000100",
INIT_01 => X"0000400000000010020311002011000000000011000203100020111800110000",
INIT_02 => X"20200000C30000000000014000000002111002001140000000010040FF000000",
INIT_03 => X"00FF18001100110000FF1800120011001400110000000000FF00022002000202",
INIT_04 => X"0000FF000003000100FF0018000011001100110000FF00180000110011001100",
INIT_05 => X"00300040002000002000D800D800FF7000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000202800000001000000",
INIT_07 => X"00000000FF00000000FF000000000000FF000000006000606000000000000000",
INIT_08 => X"00000320BE0000DE000000201100100000000010FF0000000000000000000010",
INIT_09 => X"000028000000182C000020002400002018000020000020001011003000180000",
INIT_0A => X"30000000001111002000FF1000110000000011000018FF001014FF0000000000",
INIT_0B => X"0000000000000000000000100000FF00000000000000000000FF300000002800",
INIT_0C => X"3800000000000000181100FFFF000000FF000000FFFF0000000040280011FF11",
INIT_0D => X"00000000000000000000000000FF001018100000000000000000002000000000",
INIT_0E => X"0000001000000000FF0000000010FF0000000000000000010001000000000000",
INIT_0F => X"00000000000080008803009000000000000000FF00000000001000000000FF00",
INIT_10 => X"0000000000001000008000200300000003000000000000000300000000000040",
INIT_11 => X"00000000000000200311000020031000000020031000000000888003000000FF",
INIT_12 => X"4048FF0000100000000000000010001800000000000000001000000000010020",
INIT_13 => X"00000010000000000000000000000010000010FF000038000220000000003800",
INIT_14 => X"FF00000000280000000000000010000000000000000000000000000000100000",
INIT_15 => X"020000FF00FF000300000000FF10000000000228300020000080000000000000",
INIT_16 => X"0000FF0000000010000000000300200000030000030000030000000000000080",
INIT_17 => X"000000003010101F0000000000FFFFFF00000000002030201810FF280200FF10",
INIT_18 => X"001010000000FF0000000000000020020018000000180030FFFF001000384000",
INIT_19 => X"FF000000000000800088000000FF000000000080000000FF0001000100100000",
INIT_1A => X"8088000000000000FF000000000080000000FF00000000100000800088000000",
INIT_1B => X"008800FF0000000000000000000000FF002000FF000020000000000000000000",
INIT_1C => X"2000002003110000000220000020031102002000002003110000008000000100",
INIT_1D => X"2003100000000320000020031100000020000020031102FF20000020031102FF",
INIT_1E => X"000100000000FF00000000000000001000000000400020031000000001200000",
INIT_1F => X"0140001002100000110101001002102000000000000100000001000000010000",
INIT_20 => X"01000201000201A10002010002010002014B000201000201000201651D400111",
INIT_21 => X"6C007973760000727600007300464443000D44430A4F4C204300FF1002110002",
INIT_22 => X"0000111100000069760063760072757600727576007275760072757600000D4D",
INIT_23 => X"616E616F742E424F562D756E7400727304006E00000002000000010000001111",
INIT_24 => X"000000000000000000000000000000000000000000000000757475005473612E",
INIT_25 => X"742E424F562D756E7400727304006E0000000200000001000000000000001200",
INIT_26 => X"0000000000000000000000000000000000000000757475005473612E616E616F",
INIT_27 => X"0000000000001110000000000000001000000000000000000000120000000000",
INIT_28 => X"0000000000000001121100000000000000001211000000000000000012110000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000021212",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"9C0010E800189801009800009E94009C5D94000000000000000874000008B000",
INIT_01 => X"00040018081014C05D089400009C07000908009C005D08B014009404019C0100",
INIT_02 => X"12000918500008000818D6001014009E90D05D009000EC0010E01400E8001501",
INIT_03 => X"04FD2A009000900004FD2A00A0009000A000900000000800FD000800000A000C",
INIT_04 => X"1410989C00D8004404FB042A000090009000780004FB042A0000900080007000",
INIT_05 => X"01420424012013080060125C1058FC0054504C4844403C3834302C2824201C18",
INIT_06 => X"5854504C4844403C3834302C2824201C18141000B810100004016400106400BC",
INIT_07 => X"00000001FE00000800FC020004000800FC01000400000800000801681360115C",
INIT_08 => X"00080800EF0008AD03000021A000802000080024FD0000080002000000080024",
INIT_09 => X"081C25011C1C24421C14250102141424271418250018000021A000802004011F",
INIT_0A => X"2B000800178080002403FC2528800804000480080023F47F24A3FC0000000000",
INIT_0B => X"0035000800040004000004250800E900000604000400000808F4210C1104230F",
INIT_0C => X"2100080C13001A00258000F8F4040400F3000009F8F4040400072B250D80F480",
INIT_0D => X"000800000100080C0000000800E600252525000400040004000810210008000E",
INIT_0E => X"0008002400000010EF0000080024F700000800080000000A000400FA00080002",
INIT_0F => X"040514080400251C252418251422181C240420D800000008002400000020DF00",
INIT_10 => X"280814181C202524102502252608054024000A020C0409402400060108140800",
INIT_11 => X"141C020008010425120C00082512E800030F2512D8001A000425257C1C1418E0",
INIT_12 => X"2525E80008251402010800100125092B4010FF0B000820082514181C20EC1825",
INIT_13 => X"08010C25081402000300081808001425000225F5001421014A25FF0B00002514",
INIT_14 => X"E00000080C21000C000500041021001000050008001100130013000410210200",
INIT_15 => X"9E1410E800F5013F00000000F32B001008207D25251425181C2509181C140504",
INIT_16 => X"0801FB0003000025000000182610251400260000260800260400070504000025",
INIT_17 => X"0D1A020A252326C31808001401F5FFFF01000000082A23232521FF25D814E823",
INIT_18 => X"08232BFFFF01F80109000500000025E1002100022D210525F5FF031230102101",
INIT_19 => X"E020081418081C25EC2514181CE0180810081425F31014E8007E005300250801",
INIT_1A => X"252520241014181CD8180810081425F31014E82008141825081C25EC2514181C",
INIT_1B => X"142518E0000028081014181C202400F10825ECFF010825EC0004000D00000D0A",
INIT_1C => X"000004251230013500100000062512200008000004251210040000254B08531C",
INIT_1D => X"2512DC0312000000000625125C021C0000000525125030EE00000425124020F6",
INIT_1E => X"1420181CF402E00000000020081418251C04050000042512EC04080000000006",
INIT_1F => X"040000EC20E8000094040000DC20D800000001E830201F004420040054200300",
INIT_20 => X"C00C20BB0820B8200710C00C10BB0810B8404C00C00C00BB0800B800CD00CA90",
INIT_21 => X"6C0030702F0000742F000074000D2020000A2020004E41564500FFFC5D940020",
INIT_22 => X"000080800000006F2F00302F00336E2F00326E2F00316E2F00306E2F00000A41",
INIT_23 => X"7469006400744C5245696975652E746801007500000874000008B00000008080",
INIT_24 => X"00011E0004000024A00002070B000000000000000000000074722E2E41730064",
INIT_25 => X"00744C5245696975652E746801007500000874000008B0002A00010000202000",
INIT_26 => X"04000024A00002070B000000000000000000000074722E2E4173006474690064",
INIT_27 => X"3801040000CC3C9C320130001000006CD03007012A0001000020200000011E00",
INIT_28 => X"03084D0010000010209003084800100000101080030142000100001008680308",
INIT_29 => X"00000000000000000000000000000000000000000000000053000100000020A0",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic