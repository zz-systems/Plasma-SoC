-- PLASMA_DE1_SOC.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLASMA_DE1_SOC is
	port (
		clk_clk                          : in    std_logic                     := '0';             --                       clk.clk
		hex_0_external_connection_export : out   std_logic_vector(6 downto 0);                     -- hex_0_external_connection.export
		hps_0_ddr_mem_a                  : out   std_logic_vector(14 downto 0);                    --                 hps_0_ddr.mem_a
		hps_0_ddr_mem_ba                 : out   std_logic_vector(2 downto 0);                     --                          .mem_ba
		hps_0_ddr_mem_ck                 : out   std_logic;                                        --                          .mem_ck
		hps_0_ddr_mem_ck_n               : out   std_logic;                                        --                          .mem_ck_n
		hps_0_ddr_mem_cke                : out   std_logic;                                        --                          .mem_cke
		hps_0_ddr_mem_cs_n               : out   std_logic;                                        --                          .mem_cs_n
		hps_0_ddr_mem_ras_n              : out   std_logic;                                        --                          .mem_ras_n
		hps_0_ddr_mem_cas_n              : out   std_logic;                                        --                          .mem_cas_n
		hps_0_ddr_mem_we_n               : out   std_logic;                                        --                          .mem_we_n
		hps_0_ddr_mem_reset_n            : out   std_logic;                                        --                          .mem_reset_n
		hps_0_ddr_mem_dq                 : inout std_logic_vector(31 downto 0) := (others => '0'); --                          .mem_dq
		hps_0_ddr_mem_dqs                : inout std_logic_vector(3 downto 0)  := (others => '0'); --                          .mem_dqs
		hps_0_ddr_mem_dqs_n              : inout std_logic_vector(3 downto 0)  := (others => '0'); --                          .mem_dqs_n
		hps_0_ddr_mem_odt                : out   std_logic;                                        --                          .mem_odt
		hps_0_ddr_mem_dm                 : out   std_logic_vector(3 downto 0);                     --                          .mem_dm
		hps_0_ddr_oct_rzqin              : in    std_logic                     := '0';             --                          .oct_rzqin
		plasma_soc_0_leds_ld             : out   std_logic_vector(9 downto 0);                     --         plasma_soc_0_leds.ld
		plasma_soc_0_sd_card_sd_cd       : in    std_logic                     := '0';             --      plasma_soc_0_sd_card.sd_cd
		plasma_soc_0_sd_card_sd_spi_cs   : out   std_logic;                                        --                          .sd_spi_cs
		plasma_soc_0_sd_card_sd_spi_miso : in    std_logic                     := '0';             --                          .sd_spi_miso
		plasma_soc_0_sd_card_sd_spi_mosi : out   std_logic;                                        --                          .sd_spi_mosi
		plasma_soc_0_sd_card_sd_spi_sclk : out   std_logic;                                        --                          .sd_spi_sclk
		plasma_soc_0_sd_card_sd_wp       : in    std_logic                     := '0';             --                          .sd_wp
		plasma_soc_0_switches_sw         : in    std_logic_vector(9 downto 0)  := (others => '0'); --     plasma_soc_0_switches.sw
		plasma_soc_0_uart_uart_rx        : in    std_logic                     := '0';             --         plasma_soc_0_uart.uart_rx
		plasma_soc_0_uart_uart_tx        : out   std_logic;                                        --                          .uart_tx
		sdram_controller_0_wire_addr     : out   std_logic_vector(12 downto 0);                    --   sdram_controller_0_wire.addr
		sdram_controller_0_wire_ba       : out   std_logic_vector(1 downto 0);                     --                          .ba
		sdram_controller_0_wire_cas_n    : out   std_logic;                                        --                          .cas_n
		sdram_controller_0_wire_cke      : out   std_logic;                                        --                          .cke
		sdram_controller_0_wire_cs_n     : out   std_logic;                                        --                          .cs_n
		sdram_controller_0_wire_dq       : inout std_logic_vector(15 downto 0) := (others => '0'); --                          .dq
		sdram_controller_0_wire_dqm      : out   std_logic_vector(1 downto 0);                     --                          .dqm
		sdram_controller_0_wire_ras_n    : out   std_logic;                                        --                          .ras_n
		sdram_controller_0_wire_we_n     : out   std_logic;                                        --                          .we_n
		sys_sdram_pll_0_sdram_clk_clk    : out   std_logic                                         -- sys_sdram_pll_0_sdram_clk.clk
	);
end entity PLASMA_DE1_SOC;

architecture rtl of PLASMA_DE1_SOC is
	component PLASMA_DE1_SOC_hex_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component PLASMA_DE1_SOC_hex_0;

	component PLASMA_DE1_SOC_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a       : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba      : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck      : out   std_logic;                                         -- mem_ck
			mem_ck_n    : out   std_logic;                                         -- mem_ck_n
			mem_cke     : out   std_logic;                                         -- mem_cke
			mem_cs_n    : out   std_logic;                                         -- mem_cs_n
			mem_ras_n   : out   std_logic;                                         -- mem_ras_n
			mem_cas_n   : out   std_logic;                                         -- mem_cas_n
			mem_we_n    : out   std_logic;                                         -- mem_we_n
			mem_reset_n : out   std_logic;                                         -- mem_reset_n
			mem_dq      : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs     : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n   : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt     : out   std_logic;                                         -- mem_odt
			mem_dm      : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin   : in    std_logic                      := 'X';             -- oct_rzqin
			h2f_rst_n   : out   std_logic;                                         -- reset_n
			h2f_axi_clk : in    std_logic                      := 'X';             -- clk
			h2f_AWID    : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR  : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN   : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE  : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK  : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT  : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID : out   std_logic;                                         -- awvalid
			h2f_AWREADY : in    std_logic                      := 'X';             -- awready
			h2f_WID     : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA   : out   std_logic_vector(127 downto 0);                    -- wdata
			h2f_WSTRB   : out   std_logic_vector(15 downto 0);                     -- wstrb
			h2f_WLAST   : out   std_logic;                                         -- wlast
			h2f_WVALID  : out   std_logic;                                         -- wvalid
			h2f_WREADY  : in    std_logic                      := 'X';             -- wready
			h2f_BID     : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP   : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID  : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY  : out   std_logic;                                         -- bready
			h2f_ARID    : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR  : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN   : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE  : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK  : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT  : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID : out   std_logic;                                         -- arvalid
			h2f_ARREADY : in    std_logic                      := 'X';             -- arready
			h2f_RID     : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA   : in    std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP   : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST   : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID  : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY  : out   std_logic;                                         -- rready
			f2h_axi_clk : in    std_logic                      := 'X';             -- clk
			f2h_AWID    : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR  : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN   : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE  : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK  : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT  : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY : out   std_logic;                                         -- awready
			f2h_AWUSER  : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID     : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA   : in    std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB   : in    std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST   : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID  : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY  : out   std_logic;                                         -- wready
			f2h_BID     : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP   : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID  : out   std_logic;                                         -- bvalid
			f2h_BREADY  : in    std_logic                      := 'X';             -- bready
			f2h_ARID    : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR  : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN   : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE  : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK  : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT  : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY : out   std_logic;                                         -- arready
			f2h_ARUSER  : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID     : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA   : out   std_logic_vector(127 downto 0);                    -- rdata
			f2h_RRESP   : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST   : out   std_logic;                                         -- rlast
			f2h_RVALID  : out   std_logic;                                         -- rvalid
			f2h_RREADY  : in    std_logic                      := 'X'              -- rready
		);
	end component PLASMA_DE1_SOC_hps_0;

	component plasma_soc_top is
		port (
			RST               : in  std_logic                     := 'X';             -- reset
			GCLK              : in  std_logic                     := 'X';             -- clk
			LD                : out std_logic_vector(9 downto 0);                     -- ld
			SD_CD             : in  std_logic                     := 'X';             -- sd_cd
			SD_SPI_CS         : out std_logic;                                        -- sd_spi_cs
			SD_SPI_MISO       : in  std_logic                     := 'X';             -- sd_spi_miso
			SD_SPI_MOSI       : out std_logic;                                        -- sd_spi_mosi
			SD_SPI_SCLK       : out std_logic;                                        -- sd_spi_sclk
			SD_WP             : in  std_logic                     := 'X';             -- sd_wp
			SW                : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- sw
			UART_RX           : in  std_logic                     := 'X';             -- uart_rx
			UART_TX           : out std_logic;                                        -- uart_tx
			avs_waitrequest_n : out std_logic;                                        -- waitrequest_n
			avs_response      : out std_logic_vector(1 downto 0);                     -- response
			avs_address       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			avs_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_read          : in  std_logic                     := 'X';             -- read
			avs_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_write         : in  std_logic                     := 'X';             -- write
			avs_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avm_waitrequest_n : in  std_logic                     := 'X';             -- waitrequest_n
			avm_response      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			avm_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_read          : out std_logic;                                        -- read
			avm_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_write         : out std_logic;                                        -- write
			avm_writedata     : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component plasma_soc_top;

	component PLASMA_DE1_SOC_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component PLASMA_DE1_SOC_sdram_controller_0;

	component PLASMA_DE1_SOC_sys_sdram_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component PLASMA_DE1_SOC_sys_sdram_pll_0;

	component PLASMA_DE1_SOC_mm_interconnect_0 is
		port (
			sys_sdram_pll_0_sys_clk_clk                         : in  std_logic                     := 'X';             -- clk
			plasma_soc_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			plasma_soc_0_avalon_master_0_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			plasma_soc_0_avalon_master_0_waitrequest            : out std_logic;                                        -- waitrequest
			plasma_soc_0_avalon_master_0_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			plasma_soc_0_avalon_master_0_read                   : in  std_logic                     := 'X';             -- read
			plasma_soc_0_avalon_master_0_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			plasma_soc_0_avalon_master_0_write                  : in  std_logic                     := 'X';             -- write
			plasma_soc_0_avalon_master_0_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			plasma_soc_0_avalon_master_0_response               : out std_logic_vector(1 downto 0);                     -- response
			hex_0_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			hex_0_s1_write                                      : out std_logic;                                        -- write
			hex_0_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_0_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			hex_0_s1_chipselect                                 : out std_logic;                                        -- chipselect
			sdram_controller_0_s1_address                       : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_0_s1_write                         : out std_logic;                                        -- write
			sdram_controller_0_s1_read                          : out std_logic;                                        -- read
			sdram_controller_0_s1_readdata                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_0_s1_writedata                     : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_0_s1_byteenable                    : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_0_s1_readdatavalid                 : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_0_s1_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_0_s1_chipselect                    : out std_logic                                         -- chipselect
		);
	end component PLASMA_DE1_SOC_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal sys_sdram_pll_0_sys_clk_clk                                  : std_logic;                     -- sys_sdram_pll_0:sys_clk_clk -> [hex_0:clk, hps_0:f2h_axi_clk, hps_0:h2f_axi_clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, plasma_soc_0:GCLK, rst_controller:clk, sdram_controller_0:clk]
	signal hps_0_h2f_reset_reset                                        : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal mm_interconnect_0_plasma_soc_0_avalon_master_0_waitrequest   : std_logic;                     -- mm_interconnect_0:plasma_soc_0_avalon_master_0_waitrequest -> mm_interconnect_0_plasma_soc_0_avalon_master_0_waitrequest:in
	signal plasma_soc_0_avalon_master_0_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:plasma_soc_0_avalon_master_0_readdata -> plasma_soc_0:avm_readdata
	signal plasma_soc_0_avalon_master_0_address                         : std_logic_vector(31 downto 0); -- plasma_soc_0:avm_address -> mm_interconnect_0:plasma_soc_0_avalon_master_0_address
	signal plasma_soc_0_avalon_master_0_byteenable                      : std_logic_vector(3 downto 0);  -- plasma_soc_0:avm_byteenable -> mm_interconnect_0:plasma_soc_0_avalon_master_0_byteenable
	signal plasma_soc_0_avalon_master_0_read                            : std_logic;                     -- plasma_soc_0:avm_read -> mm_interconnect_0:plasma_soc_0_avalon_master_0_read
	signal plasma_soc_0_avalon_master_0_response                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:plasma_soc_0_avalon_master_0_response -> plasma_soc_0:avm_response
	signal plasma_soc_0_avalon_master_0_write                           : std_logic;                     -- plasma_soc_0:avm_write -> mm_interconnect_0:plasma_soc_0_avalon_master_0_write
	signal plasma_soc_0_avalon_master_0_writedata                       : std_logic_vector(31 downto 0); -- plasma_soc_0:avm_writedata -> mm_interconnect_0:plasma_soc_0_avalon_master_0_writedata
	signal mm_interconnect_0_sdram_controller_0_s1_chipselect           : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	signal mm_interconnect_0_sdram_controller_0_s1_readdata             : std_logic_vector(15 downto 0); -- sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	signal mm_interconnect_0_sdram_controller_0_s1_waitrequest          : std_logic;                     -- sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_0_s1_address              : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	signal mm_interconnect_0_sdram_controller_0_s1_read                 : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_read -> mm_interconnect_0_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_0_s1_byteenable -> mm_interconnect_0_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_0_s1_readdatavalid        : std_logic;                     -- sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_0_s1_write                : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_write -> mm_interconnect_0_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_sdram_controller_0_s1_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	signal mm_interconnect_0_hex_0_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:hex_0_s1_chipselect -> hex_0:chipselect
	signal mm_interconnect_0_hex_0_s1_readdata                          : std_logic_vector(31 downto 0); -- hex_0:readdata -> mm_interconnect_0:hex_0_s1_readdata
	signal mm_interconnect_0_hex_0_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_0_s1_address -> hex_0:address
	signal mm_interconnect_0_hex_0_s1_write                             : std_logic;                     -- mm_interconnect_0:hex_0_s1_write -> mm_interconnect_0_hex_0_s1_write:in
	signal mm_interconnect_0_hex_0_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_0_s1_writedata -> hex_0:writedata
	signal rst_controller_reset_out_reset                               : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:plasma_soc_0_reset_sink_reset_bridge_in_reset_reset, plasma_soc_0:RST, rst_controller_reset_out_reset:in]
	signal sys_sdram_pll_0_reset_source_reset                           : std_logic;                     -- sys_sdram_pll_0:reset_source_reset -> rst_controller:reset_in0
	signal hps_0_h2f_reset_reset_ports_inv                              : std_logic;                     -- hps_0_h2f_reset_reset:inv -> sys_sdram_pll_0:ref_reset_reset
	signal plasma_soc_0_avalon_master_0_inv                             : std_logic;                     -- mm_interconnect_0_plasma_soc_0_avalon_master_0_waitrequest:inv -> plasma_soc_0:avm_waitrequest_n
	signal mm_interconnect_0_sdram_controller_0_s1_read_ports_inv       : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_read:inv -> sdram_controller_0:az_rd_n
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_0_s1_byteenable:inv -> sdram_controller_0:az_be_n
	signal mm_interconnect_0_sdram_controller_0_s1_write_ports_inv      : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_write:inv -> sdram_controller_0:az_wr_n
	signal mm_interconnect_0_hex_0_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_hex_0_s1_write:inv -> hex_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_reset_out_reset:inv -> [hex_0:reset_n, sdram_controller_0:reset_n]

begin

	hex_0 : component PLASMA_DE1_SOC_hex_0
		port map (
			clk        => sys_sdram_pll_0_sys_clk_clk,                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_0_s1_readdata,        --                    .readdata
			out_port   => hex_0_external_connection_export            -- external_connection.export
		);

	hps_0 : component PLASMA_DE1_SOC_hps_0
		generic map (
			F2S_Width => 3,
			S2F_Width => 3
		)
		port map (
			mem_a       => hps_0_ddr_mem_a,             --         memory.mem_a
			mem_ba      => hps_0_ddr_mem_ba,            --               .mem_ba
			mem_ck      => hps_0_ddr_mem_ck,            --               .mem_ck
			mem_ck_n    => hps_0_ddr_mem_ck_n,          --               .mem_ck_n
			mem_cke     => hps_0_ddr_mem_cke,           --               .mem_cke
			mem_cs_n    => hps_0_ddr_mem_cs_n,          --               .mem_cs_n
			mem_ras_n   => hps_0_ddr_mem_ras_n,         --               .mem_ras_n
			mem_cas_n   => hps_0_ddr_mem_cas_n,         --               .mem_cas_n
			mem_we_n    => hps_0_ddr_mem_we_n,          --               .mem_we_n
			mem_reset_n => hps_0_ddr_mem_reset_n,       --               .mem_reset_n
			mem_dq      => hps_0_ddr_mem_dq,            --               .mem_dq
			mem_dqs     => hps_0_ddr_mem_dqs,           --               .mem_dqs
			mem_dqs_n   => hps_0_ddr_mem_dqs_n,         --               .mem_dqs_n
			mem_odt     => hps_0_ddr_mem_odt,           --               .mem_odt
			mem_dm      => hps_0_ddr_mem_dm,            --               .mem_dm
			oct_rzqin   => hps_0_ddr_oct_rzqin,         --               .oct_rzqin
			h2f_rst_n   => hps_0_h2f_reset_reset,       --      h2f_reset.reset_n
			h2f_axi_clk => sys_sdram_pll_0_sys_clk_clk, --  h2f_axi_clock.clk
			h2f_AWID    => open,                        -- h2f_axi_master.awid
			h2f_AWADDR  => open,                        --               .awaddr
			h2f_AWLEN   => open,                        --               .awlen
			h2f_AWSIZE  => open,                        --               .awsize
			h2f_AWBURST => open,                        --               .awburst
			h2f_AWLOCK  => open,                        --               .awlock
			h2f_AWCACHE => open,                        --               .awcache
			h2f_AWPROT  => open,                        --               .awprot
			h2f_AWVALID => open,                        --               .awvalid
			h2f_AWREADY => open,                        --               .awready
			h2f_WID     => open,                        --               .wid
			h2f_WDATA   => open,                        --               .wdata
			h2f_WSTRB   => open,                        --               .wstrb
			h2f_WLAST   => open,                        --               .wlast
			h2f_WVALID  => open,                        --               .wvalid
			h2f_WREADY  => open,                        --               .wready
			h2f_BID     => open,                        --               .bid
			h2f_BRESP   => open,                        --               .bresp
			h2f_BVALID  => open,                        --               .bvalid
			h2f_BREADY  => open,                        --               .bready
			h2f_ARID    => open,                        --               .arid
			h2f_ARADDR  => open,                        --               .araddr
			h2f_ARLEN   => open,                        --               .arlen
			h2f_ARSIZE  => open,                        --               .arsize
			h2f_ARBURST => open,                        --               .arburst
			h2f_ARLOCK  => open,                        --               .arlock
			h2f_ARCACHE => open,                        --               .arcache
			h2f_ARPROT  => open,                        --               .arprot
			h2f_ARVALID => open,                        --               .arvalid
			h2f_ARREADY => open,                        --               .arready
			h2f_RID     => open,                        --               .rid
			h2f_RDATA   => open,                        --               .rdata
			h2f_RRESP   => open,                        --               .rresp
			h2f_RLAST   => open,                        --               .rlast
			h2f_RVALID  => open,                        --               .rvalid
			h2f_RREADY  => open,                        --               .rready
			f2h_axi_clk => sys_sdram_pll_0_sys_clk_clk, --  f2h_axi_clock.clk
			f2h_AWID    => open,                        --  f2h_axi_slave.awid
			f2h_AWADDR  => open,                        --               .awaddr
			f2h_AWLEN   => open,                        --               .awlen
			f2h_AWSIZE  => open,                        --               .awsize
			f2h_AWBURST => open,                        --               .awburst
			f2h_AWLOCK  => open,                        --               .awlock
			f2h_AWCACHE => open,                        --               .awcache
			f2h_AWPROT  => open,                        --               .awprot
			f2h_AWVALID => open,                        --               .awvalid
			f2h_AWREADY => open,                        --               .awready
			f2h_AWUSER  => open,                        --               .awuser
			f2h_WID     => open,                        --               .wid
			f2h_WDATA   => open,                        --               .wdata
			f2h_WSTRB   => open,                        --               .wstrb
			f2h_WLAST   => open,                        --               .wlast
			f2h_WVALID  => open,                        --               .wvalid
			f2h_WREADY  => open,                        --               .wready
			f2h_BID     => open,                        --               .bid
			f2h_BRESP   => open,                        --               .bresp
			f2h_BVALID  => open,                        --               .bvalid
			f2h_BREADY  => open,                        --               .bready
			f2h_ARID    => open,                        --               .arid
			f2h_ARADDR  => open,                        --               .araddr
			f2h_ARLEN   => open,                        --               .arlen
			f2h_ARSIZE  => open,                        --               .arsize
			f2h_ARBURST => open,                        --               .arburst
			f2h_ARLOCK  => open,                        --               .arlock
			f2h_ARCACHE => open,                        --               .arcache
			f2h_ARPROT  => open,                        --               .arprot
			f2h_ARVALID => open,                        --               .arvalid
			f2h_ARREADY => open,                        --               .arready
			f2h_ARUSER  => open,                        --               .aruser
			f2h_RID     => open,                        --               .rid
			f2h_RDATA   => open,                        --               .rdata
			f2h_RRESP   => open,                        --               .rresp
			f2h_RLAST   => open,                        --               .rlast
			f2h_RVALID  => open,                        --               .rvalid
			f2h_RREADY  => open                         --               .rready
		);

	plasma_soc_0 : component plasma_soc_top
		port map (
			RST               => rst_controller_reset_out_reset,          --      reset_sink.reset
			GCLK              => sys_sdram_pll_0_sys_clk_clk,             --      clock_sink.clk
			LD                => plasma_soc_0_leds_ld,                    --            leds.ld
			SD_CD             => plasma_soc_0_sd_card_sd_cd,              --         sd_card.sd_cd
			SD_SPI_CS         => plasma_soc_0_sd_card_sd_spi_cs,          --                .sd_spi_cs
			SD_SPI_MISO       => plasma_soc_0_sd_card_sd_spi_miso,        --                .sd_spi_miso
			SD_SPI_MOSI       => plasma_soc_0_sd_card_sd_spi_mosi,        --                .sd_spi_mosi
			SD_SPI_SCLK       => plasma_soc_0_sd_card_sd_spi_sclk,        --                .sd_spi_sclk
			SD_WP             => plasma_soc_0_sd_card_sd_wp,              --                .sd_wp
			SW                => plasma_soc_0_switches_sw,                --        switches.sw
			UART_RX           => plasma_soc_0_uart_uart_rx,               --            uart.uart_rx
			UART_TX           => plasma_soc_0_uart_uart_tx,               --                .uart_tx
			avs_waitrequest_n => open,                                    --  avalon_slave_0.waitrequest_n
			avs_response      => open,                                    --                .response
			avs_address       => open,                                    --                .address
			avs_byteenable    => open,                                    --                .byteenable
			avs_read          => open,                                    --                .read
			avs_readdata      => open,                                    --                .readdata
			avs_write         => open,                                    --                .write
			avs_writedata     => open,                                    --                .writedata
			avm_waitrequest_n => plasma_soc_0_avalon_master_0_inv,        -- avalon_master_0.waitrequest_n
			avm_response      => plasma_soc_0_avalon_master_0_response,   --                .response
			avm_address       => plasma_soc_0_avalon_master_0_address,    --                .address
			avm_byteenable    => plasma_soc_0_avalon_master_0_byteenable, --                .byteenable
			avm_read          => plasma_soc_0_avalon_master_0_read,       --                .read
			avm_readdata      => plasma_soc_0_avalon_master_0_readdata,   --                .readdata
			avm_write         => plasma_soc_0_avalon_master_0_write,      --                .write
			avm_writedata     => plasma_soc_0_avalon_master_0_writedata   --                .writedata
		);

	sdram_controller_0 : component PLASMA_DE1_SOC_sdram_controller_0
		port map (
			clk            => sys_sdram_pll_0_sys_clk_clk,                                  --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_0_wire_addr,                                 --  wire.export
			zs_ba          => sdram_controller_0_wire_ba,                                   --      .export
			zs_cas_n       => sdram_controller_0_wire_cas_n,                                --      .export
			zs_cke         => sdram_controller_0_wire_cke,                                  --      .export
			zs_cs_n        => sdram_controller_0_wire_cs_n,                                 --      .export
			zs_dq          => sdram_controller_0_wire_dq,                                   --      .export
			zs_dqm         => sdram_controller_0_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_controller_0_wire_ras_n,                                --      .export
			zs_we_n        => sdram_controller_0_wire_we_n                                  --      .export
		);

	sys_sdram_pll_0 : component PLASMA_DE1_SOC_sys_sdram_pll_0
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => hps_0_h2f_reset_reset_ports_inv,    --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_0_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sys_sdram_pll_0_sdram_clk_clk,      --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_0_reset_source_reset  -- reset_source.reset
		);

	mm_interconnect_0 : component PLASMA_DE1_SOC_mm_interconnect_0
		port map (
			sys_sdram_pll_0_sys_clk_clk                         => sys_sdram_pll_0_sys_clk_clk,                                --                       sys_sdram_pll_0_sys_clk.clk
			plasma_soc_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                             -- plasma_soc_0_reset_sink_reset_bridge_in_reset.reset
			plasma_soc_0_avalon_master_0_address                => plasma_soc_0_avalon_master_0_address,                       --                  plasma_soc_0_avalon_master_0.address
			plasma_soc_0_avalon_master_0_waitrequest            => mm_interconnect_0_plasma_soc_0_avalon_master_0_waitrequest, --                                              .waitrequest
			plasma_soc_0_avalon_master_0_byteenable             => plasma_soc_0_avalon_master_0_byteenable,                    --                                              .byteenable
			plasma_soc_0_avalon_master_0_read                   => plasma_soc_0_avalon_master_0_read,                          --                                              .read
			plasma_soc_0_avalon_master_0_readdata               => plasma_soc_0_avalon_master_0_readdata,                      --                                              .readdata
			plasma_soc_0_avalon_master_0_write                  => plasma_soc_0_avalon_master_0_write,                         --                                              .write
			plasma_soc_0_avalon_master_0_writedata              => plasma_soc_0_avalon_master_0_writedata,                     --                                              .writedata
			plasma_soc_0_avalon_master_0_response               => plasma_soc_0_avalon_master_0_response,                      --                                              .response
			hex_0_s1_address                                    => mm_interconnect_0_hex_0_s1_address,                         --                                      hex_0_s1.address
			hex_0_s1_write                                      => mm_interconnect_0_hex_0_s1_write,                           --                                              .write
			hex_0_s1_readdata                                   => mm_interconnect_0_hex_0_s1_readdata,                        --                                              .readdata
			hex_0_s1_writedata                                  => mm_interconnect_0_hex_0_s1_writedata,                       --                                              .writedata
			hex_0_s1_chipselect                                 => mm_interconnect_0_hex_0_s1_chipselect,                      --                                              .chipselect
			sdram_controller_0_s1_address                       => mm_interconnect_0_sdram_controller_0_s1_address,            --                         sdram_controller_0_s1.address
			sdram_controller_0_s1_write                         => mm_interconnect_0_sdram_controller_0_s1_write,              --                                              .write
			sdram_controller_0_s1_read                          => mm_interconnect_0_sdram_controller_0_s1_read,               --                                              .read
			sdram_controller_0_s1_readdata                      => mm_interconnect_0_sdram_controller_0_s1_readdata,           --                                              .readdata
			sdram_controller_0_s1_writedata                     => mm_interconnect_0_sdram_controller_0_s1_writedata,          --                                              .writedata
			sdram_controller_0_s1_byteenable                    => mm_interconnect_0_sdram_controller_0_s1_byteenable,         --                                              .byteenable
			sdram_controller_0_s1_readdatavalid                 => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,      --                                              .readdatavalid
			sdram_controller_0_s1_waitrequest                   => mm_interconnect_0_sdram_controller_0_s1_waitrequest,        --                                              .waitrequest
			sdram_controller_0_s1_chipselect                    => mm_interconnect_0_sdram_controller_0_s1_chipselect          --                                              .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_0_reset_source_reset, -- reset_in0.reset
			clk            => sys_sdram_pll_0_sys_clk_clk,        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

	plasma_soc_0_avalon_master_0_inv <= not mm_interconnect_0_plasma_soc_0_avalon_master_0_waitrequest;

	mm_interconnect_0_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_read;

	mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_write;

	mm_interconnect_0_hex_0_s1_write_ports_inv <= not mm_interconnect_0_hex_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of PLASMA_DE1_SOC
