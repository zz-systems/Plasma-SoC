---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"1000243C8C3C320CAF8C3C8CAF3C2724088C3C3C000000000003273C0003273C",
INIT_01 => X"AF24AFAF00001424AC24278C3C27038F8FA0AC242410AC240014240010240000",
INIT_02 => X"93A000932410A0009300108E3C2A020C0000001600000000001400000000AF27",
INIT_03 => X"108EA000938E00102A020C27A00093A000932410A0009300108E2A270C02A000",
INIT_04 => X"0CAF3C8E3CAF27001030008C3C00088C3C27038F8F8F8FA000838EA000838E24",
INIT_05 => X"000327083C8F8F000C8E240C3C8E240C008E240C3C8E240C008E000C8C8E3C24",
INIT_06 => X"24AC3C3CAE1000162A0C24AC24AFAE3C00243CAF248E3CAF273C14AC2C008C3C",
INIT_07 => X"243C243C241400AC243C243C241400AC243C243C273C273C0027038F8F8F2408",
INIT_08 => X"AFAFAFAFAFAF2308000C000C24142400AC8C243C243C243C24142400AC8C243C",
INIT_09 => X"8F8F8F8F8F8F8F8F8F8F8F000CAF00AF00AF2340AFAFAFAFAFAFAFAFAFAFAFAF",
INIT_0A => X"001030008C0003001030008C0040034040033423038F038F8F8F8F8F8F8F8F8F",
INIT_0B => X"AFAFAFAFAF3CAF270003AC00248C0003AC34008C0003AC00008CAC34248C0003",
INIT_0C => X"8F8F8F2616263C0C0202000010008E00120014020210028E24243C000026AFAF",
INIT_0D => X"8F028F8F003C0C3002003C0C02AC0024AFAF00240030AF3C2727038F8F8F8F8F",
INIT_0E => X"00008C0010248C3C0024240010AC03ACACAC24AC3C00343C0024243C27083C30",
INIT_0F => X"3C100003ACACACAC008C8C000300108CAC10ACACAC008CACAC240024142C0014",
INIT_10 => X"00008C241000108C008CACACACAC8C00108CAC10ACACAC8C001100001024248C",
INIT_11 => X"00248C000300248C0000000300108C000000ACACACAC008C8CAC2400008C0014",
INIT_12 => X"AC0000308CAC0000008C240003AC0000308CAC0000008C240003AC00008CAC00",
INIT_13 => X"AC00248C0003AC340003ACAC340003AC000003AC0000308CAC0000008C240003",
INIT_14 => X"0003AC34008C000800080008000003AC0003AC00341024108C0003AC0000308C",
INIT_15 => X"AF8CAF2700000003AC00008CAC34248C0003AC00008CAC34248C0003AC00248C",
INIT_16 => X"24AEAE243C16240010AEAE24AEAE243C1624ACACACAC0010000C2400AF12AFAF",
INIT_17 => X"24AE10240C0012001232AEAE240010020CAE14240C00100010322424001024AE",
INIT_18 => X"3C10020C243C2410020C243C10008C00000CAFAFAF2727038F8F8F8F028FAEAE",
INIT_19 => X"AC24001000008C8C3010008C2703008F8F8F27088F028F8F2400102410020C24",
INIT_1A => X"2703008F0000100010008D00250C013010008100AF000027000300AC242403A0",
INIT_1B => X"100014008CAC0010008C2414000300AC24000390AC24001000008C8C0010008C",
INIT_1C => X"10008CAC0000008C0010008C001400108C0010008CAC00008C0010008C241400",
INIT_1D => X"8E001002008E8C270800008F028F8F0014AFAFAF248C278C0003AC0000008C00",
INIT_1E => X"0027088F028F000C8E000C8E000C8E0010248C008E000CAFAF270010260C8C92",
INIT_1F => X"2703008FA01024A02480800010000000000024000CAF27000324100010008000",
INIT_20 => X"1000140080800008A000A1242400040010A11000240000240000152400000000",
INIT_21 => X"8F8E8F000CAFAF27000800080003A01424802400000003340300003030241024",
INIT_22 => X"AFAF2727038F8F00AE8F000C00AFAFAF2727038F8FAE8F000C00AFAFAF272703",
INIT_23 => X"AE020C8226AE020C00140010008224240000AFAFAFAFAFAF2727038F8E8F000C",
INIT_24 => X"24103C3C14020C24ACAC3C0010240CAFAF00AF27000027038F8F8F8F8F8F0010",
INIT_25 => X"3C3C14020C2424103C3C14020C2424103C3C14020C242410AE243C3C14020C24",
INIT_26 => X"8FAE24AE3C14020C242410AE243C3C14020C242410AE243C3C14020C242410AE",
INIT_27 => X"240C243C240C243C240C243C240C243CAF0CAFAF2400273C00000027038F8F02",
INIT_28 => X"3C3C0C3C0C3C0CAC0C3C3C240C243C3CAE0C263C240C243C3C3C240C240C243C",
INIT_29 => X"260C24360C24360C24260C343C360C24360C24260C243C360C24360C24260C24",
INIT_2A => X"77307564724F4C494F4C493A5421544953410010240C8E3C360C360C24360C24",
INIT_2B => X"64006964007463640074636400746364007463647200303000496F48006C6464",
INIT_2C => X"00000F410003273C0003273C0000000000000000000000000000000000003067",
INIT_2D => X"000000000000006569616743002E6161742E612E65455443646C2E2E6E617300",
INIT_2E => X"65455443646C2E2E6E61730000000F410003273C0003273C0000000000000000",
INIT_2F => X"000000000000000000000000000000000000006569616743002E6161742E612E",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"4062420283040500BF440250B002BDA5004405020000000000405A1A00405A1A",
INIT_01 => X"B112B2B0074360036242BD6203BDE0B0BF6285650200A2620046068046060210",
INIT_02 => X"A34300A303004300A3006002100300000007524000000007836000000000BFA5",
INIT_03 => X"00024300A3020040424000A54300A34300A303004300A300800224A500204300",
INIT_04 => X"00BF050410B0BD00404200420200004402BDE0B0B1B2BF4300A3024300A30203",
INIT_05 => X"00E0BD0004B0BF000004A500050405000004A5000504050000040000450402A5",
INIT_06 => X"A54005022000000010008443A5BF3002627005B0022311B1BD04406444006203",
INIT_07 => X"A505C606A560A4A08404A505A560A4A08404A505BD1D9C1C00BDE0B0B1BF8400",
INIT_08 => X"A6A5A4A3A2A1BD0000000000A560C6A4A3C38404A505C606A560C6A4A3C38404",
INIT_09 => X"ABAAA9A8A7A6A5A4A3A2A10000BB00BB00BA5A1ABFB9B8AFAEADACABAAA9A8A7",
INIT_0A => X"004042008200E000404200820084E0029B401BBD60BB60BBBABFB9B8AFAEADAC",
INIT_0B => X"B0B3B4B5B611B1BD00E08243038200E08242008200E0824300828242038200E0",
INIT_0C => X"B5B6BF3114100400007240004000220040004053424016A2141615000031B2BF",
INIT_0D => X"B120B0BF100400C6201004002044A006B0BF624211B1B102BDBDE0B0B1B2B3B4",
INIT_0E => X"A400650062424302828402008082E043436283430462630343420302BD0004C6",
INIT_0F => X"038000E0606085A400656400E00000636600C3C486006464C5A54462C0A6A4C0",
INIT_10 => X"E4006467600045460062468287E6E2000042E600878246470000C2E047678662",
INIT_11 => X"A20283A2E0A30382000000E00000C6C04060404087E400444764848700470047",
INIT_12 => X"85A2A6C682824302A2830200E085A2A6C682824302A2830200E085A2058283A3",
INIT_13 => X"8243038200E085A500E08582A200E0850000E085A2A6C682824302A2830200E0",
INIT_14 => X"00E0824200820000000000000000E08500E08243420003A08200E085A205A582",
INIT_15 => X"BF93B3BD000000E0824300828242038200E0824300828242038200E082430382",
INIT_16 => X"020202420262020000000202020242026202404040524040A0000480B060B1B2",
INIT_17 => X"0302400400004000203102030300000000024004000040006023021200001202",
INIT_18 => X"05400000A50505400000A50540004240A000BFB0B1BDBDE0B0B1B2B300BF0203",
INIT_19 => X"82C20060C2438683A5400082BDE000B0B1BFBD00B120B0BF05000005400000A5",
INIT_1A => X"BDE000BF000000E0400022E2080020A5A0000500BFA080BD00E000820202E0C5",
INIT_1B => X"0000400082824540008202C000E000820200E0A282A20060A243858300400082",
INIT_1C => X"4000828243A300830040008200C245008200400082824500820040008202C200",
INIT_1D => X"02004022000291BD000000B000B1BF8062B1BFB00243BD8200E08545A3008300",
INIT_1E => X"00BD00B000BF0000040000040000040062024300028000BFB0BD000031004425",
INIT_1F => X"BDE000BF4400426663466400808645658082428000BFBD44E042000060004380",
INIT_20 => X"40004300A382A00060A302C302A3816000074000E700A3C30749200900436404",
INIT_21 => X"B002BF8000B0BFBD0000000000E0648063A4A5808000E042E002434263A50084",
INIT_22 => X"B0BFBDBDE0B0B10011BF8000A0B0B1BFBDBDE0B0B111BF8000A0B0B1BFBDBDE0",
INIT_23 => X"34200014103320000052004000021312A080B4BFB0B1B2B3BDBDE0B002BF8000",
INIT_24 => X"42000205402000A540400540400400BFB080B1BD0000BDE0B0B1B2B3B4BF0000",
INIT_25 => X"0205402000A542000205402000A542000205402000A5020002420205402000A5",
INIT_26 => X"BF02020202402000A5020002420205402000A5020002420205402000A5020002",
INIT_27 => X"84000504840005048400050484000504B000B1BF8400BD04000000BDE0B0B100",
INIT_28 => X"05040004000400620004038400A50405220004118400A5100405040084000504",
INIT_29 => X"0400050400050400050400A5050400050400050400A5050400050400050400A5",
INIT_2A => X"00006165774645524E455220690D494F53430000A50024050400040005040005",
INIT_2B => X"6500726500656F6500656F6500656F6500656F6500003A30004E206500616965",
INIT_2C => X"0701670000405A1A00405A1A0000000000000000000000000000000000000070",
INIT_2D => X"000000000000007362746E4B536274006469747278004154006462676F62742E",
INIT_2E => X"78004154006462676F62742E0701670000405A1A00405A1A0000000000000000",
INIT_2F => X"000000000000000000000000000000000000007362746E4B5362740064697472",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"0010160016000003001600010020FF1503160000000000000000040000000300",
INIT_01 => X"000E0000000000001600FF160000000000001600000016FF0000002800001616",
INIT_02 => X"0000000000000000000000160000200490000000000088000000000080200000",
INIT_03 => X"0016000000160000002004000000000000000000000000000016000004200000",
INIT_04 => X"030000160000FF00000000004000031600000000000000000000160000001600",
INIT_05 => X"0000000240000000031616030016000330161603001600033016000316160015",
INIT_06 => X"150400201600000000041604150016201800000000160000FF00001600001600",
INIT_07 => X"1600160000FF18001600160000FF180017001600190016000000000000001604",
INIT_08 => X"000000000000FF010004000100FF0018000016001600160000FF001800001600",
INIT_09 => X"0000000000000000000000000100D800D800FF70000000000000000000000000",
INIT_0A => X"00FF000000000000FF0000000060006060000000000000000000000000000000",
INIT_0B => X"00000000000000FF00000010FF000000000000000000001000000000FF000000",
INIT_0C => X"00000000FF0020022898F8000000000000000010900090000000209880160000",
INIT_0D => X"002800003420020028342002280080000000101618000000FF00000000000000",
INIT_0E => X"30000000001616002000FF1000160000000016000018FF001019FF0000022000",
INIT_0F => X"0000000000000000000000100000FF00000000000000000000FF300000002800",
INIT_10 => X"3800000000000000181600FFFF000000FF000000FFFF0000000040280016FF16",
INIT_11 => X"28000010002800000000000000FF001018100000000000000000002000000000",
INIT_12 => X"0028280000001010100000000000282800000010101000000000002828000018",
INIT_13 => X"0010FF0000000000000000000000000000000000282800000010101000000000",
INIT_14 => X"00000000000000010001000100000000000000100000FF000000000028280000",
INIT_15 => X"000000FF00000000001000000000FF000000001000000000FF0000000010FF00",
INIT_16 => X"0000000120000090000000000000004000000000000080008804009000000000",
INIT_17 => X"0000FF0004000000000000000080002004000000040000000000000010000000",
INIT_18 => X"000020041500000020041500000000888004000000FF00000000000010000000",
INIT_19 => X"0000100018100000000000000000100000000002002000000000000000200415",
INIT_1A => X"0000000010000010FF0000380003200000000038004048FF0000100000000000",
INIT_1B => X"0000000000001000000000000000100000000000000010001810000000000000",
INIT_1C => X"0000000010180000000000000000280000000000000010000000000000000000",
INIT_1D => X"0000FF10000000000328300020000080000000000000FF000000002828000000",
INIT_1E => X"00000400200000040000040000040000000000000080030000FF00FF00040000",
INIT_1F => X"0000000000FFFFFF00000000002030201810FF280300FF100000FF0000000010",
INIT_20 => X"00000000000020030018000000180030FFFF001000384000000000003010101F",
INIT_21 => X"00000080010000FF000100010000FFFF00FF001810100000001010000000FF00",
INIT_22 => X"0000FF00000000100000800188000000FF000000000000800188000000FF0000",
INIT_23 => X"002001FF0000200100000000000000008088000000000000FF00000000008001",
INIT_24 => X"03002000002004150000008000000100008800FF0000000000000000000000FF",
INIT_25 => X"20000020041503FF20000020041503FF20000020041500000003200000200415",
INIT_26 => X"0000000040002004150000000120000020041500000004200000200415000000",
INIT_27 => X"02010000030100000201000000010000000100000028FF000000000000000010",
INIT_28 => X"0040014002400216014000150315000016010100150315200000000100010000",
INIT_29 => X"0202000302000302000302A10003020003020003025E00030200030200030212",
INIT_2A => X"0000727600464443204443006D0A4F4C204300FF150316000201020203020200",
INIT_2B => X"76006376007275760072757600727576007275760000303A000D4D6C00797376",
INIT_2C => X"04006E0000000400000003000000161600001516000016160000151600000069",
INIT_2D => X"0000000000000000757475005473612E616E616F742E424F562D756E74007273",
INIT_2E => X"742E424F562D756E7400727304006E0000000400000003000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000757475005473612E616E616F",
INIT_30 => X"0000000000001515000000000000001500000000000000000000160000000000",
INIT_31 => X"0000000000000000161600000000000000001616000000000000000016160000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000021617",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"0F2B70003000FF34148400081000E8384884000000000000000864000008A000",
INIT_01 => X"1C1020180D1A023C8801D8880018081014003001200330FF00057F2504080300",
INIT_02 => X"100700113006070010000634000A2500120D1A020000100D1A02000010122410",
INIT_03 => X"08340100103400080A25001003001004001130060400100006340A1000250600",
INIT_04 => X"481400800010E800260100040000A884002808181C2024000010340100113430",
INIT_05 => X"000818A600101400A8805048008020742580704800801074258000483480004C",
INIT_06 => X"6008000090070009082B7008541C90000401001401900018E000168C01008C00",
INIT_07 => X"3000100004FD2A005000500004FD2A00200050002000500000200814181C702B",
INIT_08 => X"24201C181410981800E800C404FB042A000050005000280004FB042A00005000",
INIT_09 => X"3834302C2824201C181410007860125C1058FC0054504C4844403C3834302C28",
INIT_0A => X"00FC020004000800FC01000400000800000801681360115C5854504C4844403C",
INIT_0B => X"101C2024280014D000080024FD000008000200000008002400000001FE000008",
INIT_0C => X"24282C04EC01003D25250900060000000A000C24241204082001002525A0182C",
INIT_0D => X"1825141C420055012502004825002501141C21A0801F1800E030081014181C20",
INIT_0E => X"2B000800174040002403FC2528400804000440080023F47F2423FC0020620001",
INIT_0F => X"0035000800040004000004250800E900000604000400000808F4210C1104230F",
INIT_10 => X"2100080C13001A00254000F8F4040400F3000009F8F4040400072B250D40F440",
INIT_11 => X"04011024080401000000000800E600252525000400040004000810210008000E",
INIT_12 => X"1425040114142427041401000818250401181824270418010008102427101025",
INIT_13 => X"0024C70000080002000800000100080C0000081C2504011C1C2427041C010008",
INIT_14 => X"0008000800000072006C00620000080C000800240402FB030000080025C00700",
INIT_15 => X"240420D800000008002400000020DF000008002400000010EF0000080024F700",
INIT_16 => X"010C0408000905250A1418401008080009061C080400252825342025142E181C",
INIT_17 => X"4008F140340008000A020C14402510253604054034000C000E01010125030114",
INIT_18 => X"0008251A7C00030F251A6C001A000425258C1C1418E0280814181C2025241018",
INIT_19 => X"100125092B211018FF0C000820082514181C20BC1825141C0200080104251AAC",
INIT_1A => X"1808001425000225F5001C21013425FF0B000025142525E80008251C02010800",
INIT_1B => X"26002600041021020008010C0008251C020008000C0125042B210C14000C0004",
INIT_1C => X"060004102121001800060008001321140C001800041021001000050008021000",
INIT_1D => X"0000F32B001008207425251425181C2509181C140604E00000080C2121001400",
INIT_1E => X"00183610251400360000360800360400070604000025A81410E800F5014F0000",
INIT_1F => X"1808001401F5FFFF01000000082A23232521FF25E014E8230801FB0003000025",
INIT_20 => X"09000500000025E9002100022D210525F5FF0312301021010D1A020A252326C3",
INIT_21 => X"100814255B1014E800FE00D30008FFFC01FF01252525080108232BFFFF01F801",
INIT_22 => X"1014E82008141825081C25542514181CE020081418081C25542514181CE01808",
INIT_23 => X"082554FF010825540004000D00000D0A252520241014181CD81808100814255B",
INIT_24 => X"0008000004251AB0040000254B08D31C142518E0000028081014181C202400F1",
INIT_25 => X"000005251AF030EE000004251AE020F6000004251AD001350010000006251AC0",
INIT_26 => X"1C0406000004251A8005080000000006251A7004120000000006251AFC031C00",
INIT_27 => X"3CA7080000A707004CA70600CCA7020014A7181C4425E0000000002008141825",
INIT_28 => X"13005400B0009A806C0000800A7C0000846C0000700A6C000000015030A71F00",
INIT_29 => X"007C0320780C2073082070200710780C1073081070105F00780C0073080070D0",
INIT_2A => X"0000742F000020200020200065004E41564500FF90488400006C0090E8008701",
INIT_2B => X"2F00302F00336E2F00326E2F00316E2F00306E2F00003030000A416C0030702F",
INIT_2C => X"01007500000864000008A000000040400000A050000040400000A0500000006F",
INIT_2D => X"000000000000000074722E2E417300647469006400744C5245696975652E7468",
INIT_2E => X"00744C5245696975652E746801007500000864000008A000A00002070B000000",
INIT_2F => X"04000024A00002070B000000000000000000000074722E2E4173006474690064",
INIT_30 => X"3801040000D0D8383201300010000008D03007012A0001000020D00000011E00",
INIT_31 => X"03084D00100000D0D0500308480010000020B0300301420001000020A8080308",
INIT_32 => X"000000000000000000000000000000000000000000000000530001000000D020",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic