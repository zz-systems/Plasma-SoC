---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"8E3CAF273C14AC2C008C3C00088C3C24088C3C3C000000000003273C0003273C",
INIT_01 => X"3CAF3C2727038F8F8F240824AC3C3CAE1000162A0C24AC24AFAE3C00243CAF24",
INIT_02 => X"1002008E00162402122400300C008C3C001402263CAF14AFAFAFAF00243C8E8C",
INIT_03 => X"3C8E3CAF27001030008C3C27038F8F8F8F8F8FA0AE241200008EA01024AC243C",
INIT_04 => X"27083C8F8F000C8E240C3C8E240C008E240C3C8E240C008E000C8C8E3C240CAF",
INIT_05 => X"AF8CAF3C2727038FA28F8FA200932410A20012932A0CAF020027AF00AF270003",
INIT_06 => X"8F8E8F8F8F8F00021424240C000002168EAC0C0000AF24AF8E3CAF0002162426",
INIT_07 => X"AC8C243C243C243C241400AC243C243C241400AC243C243C273C273C00270800",
INIT_08 => X"AFAFAFAFAFAFAFAFAFAF2308000C000C24142400AC8C243C243C243C24142400",
INIT_09 => X"8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F000CAF00AF00AF2340AFAFAFAFAFAFAFAF",
INIT_0A => X"248C0003001030008C0003001030008C0040034040033423038F038F8F8F8F8F",
INIT_0B => X"ACAC3C0010240CAFAF00AF270003AC00248C0003AC34008C0003AC00008CAC34",
INIT_0C => X"3C14020C2424103C3C14020C24AE1024AE243C3C14020C2424103C3C14020C24",
INIT_0D => X"2410AE243C3C14020C242410AE243C3C14020C242410AE3C3C14020C2424103C",
INIT_0E => X"AF3CAF2700000010000CAF2700000027038F8F028F00020C2410AE3C14020C24",
INIT_0F => X"16263C0C0202000010008E00120014020210028E24243C000026AFAFAFAFAFAF",
INIT_10 => X"003C0C3002003C0C02AC0024AFAF00240030AF3C2727038F8F8F8F8F8F8F8F26",
INIT_11 => X"10248C3C0024240010AC03ACACAC24AC3C00343C0024243C27083C308F028F8F",
INIT_12 => X"ACACACAC008C8C000300108CAC10ACACAC008CACAC240024142C001400008C00",
INIT_13 => X"1000108C008CACACACAC8C00108CAC10ACACAC8C001100001024248C3C100003",
INIT_14 => X"0300248C0000000300108C000000ACACACAC008C8CAC2400008C001400008C24",
INIT_15 => X"8CAC0000008C240003AC0000308CAC0000008C240003AC00008CAC0000248C00",
INIT_16 => X"0003AC340003ACAC340003AC000003AC0000308CAC0000008C240003AC000030",
INIT_17 => X"008C000800080008000003AC0003AC00341024108C0003AC0000308CAC00248C",
INIT_18 => X"00000003AC00008CAC34248C0003AC00008CAC34248C0003AC00248C0003AC34",
INIT_19 => X"3C16240010AEAE24AEAE243C1624ACACACAC0010000C2400AF12AFAFAF8CAF27",
INIT_1A => X"0C0012001232AEAE240010020CAE14240C00100010322424001024AE24AEAE24",
INIT_1B => X"243C2410020C243C10008C00000CAFAFAF2727038F8F8F8F028FAEAE24AE1024",
INIT_1C => X"00008C8C3010008C2703008F8F8F27088F028F8F2400102410020C243C10020C",
INIT_1D => X"0000100010008D00250C013010008100AF000027000300AC242403A0AC240010",
INIT_1E => X"8CAC0010008C2414000300AC24000390AC24001000008C8C0010008C2703008F",
INIT_1F => X"0000008C0010008C001400108C0010008CAC00008C0010008C24140010001400",
INIT_20 => X"008E8C270800008F028F8F0014AFAFAF248C278C0003AC0000008C0010008CAC",
INIT_21 => X"028F000C8E000C8E000C8E0010248C008E000CAFAF270010260C8C928E001002",
INIT_22 => X"A01024A02480800010000000000024000CAF270003241000100080000027088F",
INIT_23 => X"80800008A000A1242400040010A110002400002400001524000000002703008F",
INIT_24 => X"0CAFAF27000800080003A0142480240000000334030000303024102410001400",
INIT_25 => X"038F8F00AE8F000C30AFAFAF2727038F8FAE8F000C00AFAFAF2727038F8E8F00",
INIT_26 => X"AE020C00140010008224240000AFAFAFAFAFAF272703308F8F8E000CAFAF2727",
INIT_27 => X"240C243C240C243CAF0CAFAF2400273C0027038F8F8F8F8F8F0010AE020C9226",
INIT_28 => X"0C3C3C240C243C3CAE0C263C240C243C3C3C240C240C243C240C243C240C243C",
INIT_29 => X"36340C263C240C36240C36240C263C240C36240C36240C263C3C0C3C0C3C0CAC",
INIT_2A => X"8F8F240C243C3C240C3C8C3C240C3C8E360C360C24240C36240C26240C36240C",
INIT_2B => X"30300D4D6C0D006C646477307564723A544F4C494F4C4921544953412703008F",
INIT_2C => X"0000000000000000723067640069640074636400746364007463640074636400",
INIT_2D => X"65455443646C2E2E6E61730000000F410003273C0003273C0000000000000000",
INIT_2E => X"0003273C0000000000000000000000000000006569616743002E6161742E612E",
INIT_2F => X"69616743002E6161742E612E65455443646C2E2E6E61730000000F410003273C",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000065",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"2311B1BD0440644400620300004402A5004405020000000000405A1A00405A1A",
INIT_01 => X"12B202BDBDE0B0B1BF8400A54005022000000010008443A5BF3002627005B002",
INIT_02 => X"4003008300620240620213A5000544024060233111B080B1B3B4BF6242024345",
INIT_03 => X"050410B0BD004042004202BDE0B0B1B2B3B4BF53434320510042620002446402",
INIT_04 => X"BD0004B0BF000004A500050405000004A5000504050000040000450402A500BF",
INIT_05 => X"B150B002BDBDE0B002B1BF0300A30200020020A23100BF2080A5B0A0B1BD00E0",
INIT_06 => X"B244B0B1B3BF0705A0058400000771204450000000BF84B34412B20711201110",
INIT_07 => X"A3C38404A505C606A560A4A08404A505A560A4A08404A505BD1D9C1C00BD0000",
INIT_08 => X"AAA9A8A7A6A5A4A3A2A1BD0000000000A560C6A4A3C38404A505C606A560C6A4",
INIT_09 => X"AFAEADACABAAA9A8A7A6A5A4A3A2A10000BB00BB00BA5A1ABFB9B8AFAEADACAB",
INIT_0A => X"038200E0004042008200E000404200820084E0029B401BBD60BB60BBBABFB9B8",
INIT_0B => X"40400540400400BFB080B1BD00E08243038200E08242008200E0824300828242",
INIT_0C => X"05402000A542000205402000A502000202420205402000A542000205402000A5",
INIT_0D => X"020002420205402000A5020002420205402000A50200020205402000A5420002",
INIT_0E => X"B611B1BD000000000000BFBD000000BDE0B0B100BF00000002000202402000A5",
INIT_0F => X"14100400007240004000220040004053424016A2141615000031B2BFB0B3B4B5",
INIT_10 => X"100400C6201004002044A006B0BF624211B1B102BDBDE0B0B1B2B3B4B5B6BF31",
INIT_11 => X"62424302828402008082E043436283430462630343420302BD0004C6B120B0BF",
INIT_12 => X"606085A400656400E00000636600C3C486006464C5A54462C0A6A4C0A4006500",
INIT_13 => X"600045460062468287E6E2000042E600878246470000C2E047678662038000E0",
INIT_14 => X"E0A30382000000E00000C6C04060404087E400444764848700470047E4006467",
INIT_15 => X"82824302A2830200E085A2A6C682824302A2830200E085A2058283A3A20283A2",
INIT_16 => X"00E085A500E08582A200E0850000E085A2A6C682824302A2830200E085A2A6C6",
INIT_17 => X"00820000000000000000E08500E08243420003A08200E085A205A58282430382",
INIT_18 => X"000000E0824300828242038200E0824300828242038200E08243038200E08242",
INIT_19 => X"0262020000000202020242026202404040524040A0000480B060B1B2BF93B3BD",
INIT_1A => X"0000400020310203030000000002400400004000602302120000120202020242",
INIT_1B => X"A50505400000A50540004240A000BFB0B1BDBDE0B0B1B2B300BF020303024004",
INIT_1C => X"C2438683A5400082BDE000B0B1BFBD00B120B0BF05000005400000A505400000",
INIT_1D => X"000000E0400022E2080020A5A0000500BFA080BD00E000820202E0C582C20060",
INIT_1E => X"82824540008202C000E000820200E0A282A20060A243858300400082BDE000BF",
INIT_1F => X"43A300830040008200C245008200400082824500820040008202C20000004000",
INIT_20 => X"000291BD000000B000B1BF8062B1BFB00243BD8200E08545A300830040008282",
INIT_21 => X"00BF0000040000040000040062024300028000BFB0BD00003100442502004022",
INIT_22 => X"4400426663466400808645658082428000BFBD44E04200006000438000BD00B0",
INIT_23 => X"A382A00060A302C302A3816000074000E700A3C30749200900436404BDE000BF",
INIT_24 => X"00B0BFBD0000000000E0648063A4A5808000E042E002434263A5008440004300",
INIT_25 => X"E0B0B10011BF8000B1B0B1BFBDBDE0B0B111BF8000A0B0B1BFBDBDE0B002BF80",
INIT_26 => X"3320000052004000021312A080B4BFB0B1B2B3BDBDE042B0BF028000BFB0BDBD",
INIT_27 => X"8400050484000504B000B1BF8400BD0400BDE0B0B1B2B3B4BF00003420001410",
INIT_28 => X"0004038400A50405220004118400A51004050400840005048400050484000504",
INIT_29 => X"04A5000405050004050004A5000405050004050004A500040504000400040062",
INIT_2A => X"B1BF8400A50405A500054402A500052404000400050500040500040500040500",
INIT_2B => X"3A300A416C0A00616965000061657720694645524E45520D494F5343BDE000B0",
INIT_2C => X"00000000000000000000706500726500656F6500656F6500656F6500656F6500",
INIT_2D => X"78004154006462676F62742E0701670000405A1A00405A1A0000000000000000",
INIT_2E => X"00405A1A0000000000000000000000000000007362746E4B5362740064697472",
INIT_2F => X"62746E4B536274006469747278004154006462676F62742E0701670000405A1A",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000073",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"160000FF00001600001600000416001503160000000000000000040000000300",
INIT_01 => X"000020FF00000000001604150400201600000000041604150016201800000000",
INIT_02 => X"00100016000000A000009E00039E160080001816000000000000002016001601",
INIT_03 => X"00160000FF000000000040000000000000000000160000880016FF000016FF00",
INIT_04 => X"0003400000000416160300160003301616030016000330160003161600150300",
INIT_05 => X"00160000FF000000000000000000000000000000000400208000008800FF0000",
INIT_06 => X"0016000000000000000E00002800000016160098280000001600000000000000",
INIT_07 => X"000016001600160000FF18001600160000FF1800170016001900160000000028",
INIT_08 => X"00000000000000000000FF010001000200FF0018000016001600160000FF0018",
INIT_09 => X"000000000000000000000000000000000100D800D800FF700000000000000000",
INIT_0A => X"FF00000000FF000000000000FF00000000600060600000000000000000000000",
INIT_0B => X"0000008000000200008800FF00000010FF000000000000000000001000000000",
INIT_0C => X"000020041603FF20000020041600000000032000002004160300200000200416",
INIT_0D => X"00FF000120000020041500FF000420000020041600FF0020000020041603FF20",
INIT_0E => X"000000FF000000FF000400FF00000000000000100080200200FF004000200415",
INIT_0F => X"FF0020022898F800000000000000001090009000000020988016000000000000",
INIT_10 => X"3420020028342002280080000000101618000000FF0000000000000000000000",
INIT_11 => X"001616002000FF1000160000000016000018FF001019FF000002200000280000",
INIT_12 => X"00000000000000100000FF00000000000000000000FF30000000280030000000",
INIT_13 => X"00000000181600FFFF000000FF000000FFFF0000000040280016FF1600000000",
INIT_14 => X"002800000000000000FF00101810000000000000000000200000000038000000",
INIT_15 => X"0000101010000000000028280000001010100000000000282800001828000010",
INIT_16 => X"0000000000000000000000000000000028280000001010100000000000282800",
INIT_17 => X"000000010001000100000000000000100000FF0000000000282800000010FF00",
INIT_18 => X"00000000001000000000FF000000001000000000FF0000000010FF0000000000",
INIT_19 => X"20000090000000000000004000000000000080008804009000000000000000FF",
INIT_1A => X"0400000000000000008000200400000004000000000000001000000000000001",
INIT_1B => X"1500000020041500000000888001000000FF000000000000100000000000FF00",
INIT_1C => X"1810000000000000000010000000000300200000000000000020041600002004",
INIT_1D => X"10000010FF0000380003200000000038004048FF000010000000000000001000",
INIT_1E => X"0000100000000000000010000000000000001000181000000000000000000000",
INIT_1F => X"1018000000000000000028000000000000001000000000000000000000000000",
INIT_20 => X"000000000328300020000080000000000000FF00000000282800000000000000",
INIT_21 => X"200000040000040000040000000000000080040000FF00FF000400000000FF10",
INIT_22 => X"00FFFFFF00000000002030201810FF280400FF100000FF000000001000000400",
INIT_23 => X"000020040018000000180030FFFF001000384000000000003010101F00000000",
INIT_24 => X"010000FF000200020000FFFF00FF001810100000001010000000FF0000000000",
INIT_25 => X"000000100000800100000000FF000000000000800188000000FF000000000080",
INIT_26 => X"00200100000000000000008088000000000000FF00000000000080010000FF00",
INIT_27 => X"0102000002020000000200000028FF0000000000000000000000FF002001FF00",
INIT_28 => X"0140001503150000160101001503152000000001000200000002000000020000",
INIT_29 => X"03A10203000002030002035E0203000002030002031202030040014003400216",
INIT_2A => X"0000160416000015040016001503001602010202000002020002020002030002",
INIT_2B => X"303A00496F48007973760000727600006D4644432044430A4F4C204300001000",
INIT_2C => X"0000161600001516000069760063760072757600727576007275760072757600",
INIT_2D => X"742E424F562D756E7400727304006E0000000400000003000000161600001516",
INIT_2E => X"0000030000000000000000000000000000000000757475005473612E616E616F",
INIT_2F => X"757475005473612E616E616F742E424F562D756E7400727304006E0000000400",
INIT_30 => X"0000000000001700000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000171600000000000000001615000000000000001500000000",
INIT_32 => X"0000000000000000000217170000000000000000171600000000000000001716",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"E00018E00016DC0100DC00000CD40090ACD40000000000000008540000089000",
INIT_01 => X"001800D8200814181CC08FB0080000E0070009088FC008A41CE0000401001401",
INIT_02 => X"0D2B0080000B7F25040803FF9800D400251E2BC0001023141C20242BA0008008",
INIT_03 => X"00D00010E800260100040028081014181C2024008001032B0080FF082080FF00",
INIT_04 => X"180A001014000CD0A0AC00D020D825D0C0AC00D010D825D000AC84D000BCAC14",
INIT_05 => X"18D81400D828081C0020240100113004010004100A64242525101C2520D80008",
INIT_06 => X"1C84141820240D1A021003A2100D1A0284D8A2121024062084001C0D1A023C01",
INIT_07 => X"0000A0008000600004FD2A00A000A00004FD2A007000A0007000A0000028A212",
INIT_08 => X"34302C2824201C181410981400D4002804FB042A0000A000A000800004FB042A",
INIT_09 => X"4844403C3834302C2824201C18141000DC60125C1058FC0054504C4844403C38",
INIT_0A => X"FE00000800FC020004000800FC01000400000800000801681360115C5854504C",
INIT_0B => X"040000254F08371C142518E000080024FD000008000200000008002400000001",
INIT_0C => X"0004257E3420F5000004257E240439010010000007257E140008000004257E04",
INIT_0D => X"05D20000000006257EC804DC0000000006257E5003E600000005257E4430ED00",
INIT_0E => X"280014D0000000FF00F014E800000020081418251C25256207CA000004257ED8",
INIT_0F => X"EC0100A125250900060000000A000C24241204082001002525F0182C101C2024",
INIT_10 => X"4200B901250200AC25002501141C21F0801F1800E030081014181C2024282C04",
INIT_11 => X"179090002403FC2528900804000490080023F47F2473FC0020C600011825141C",
INIT_12 => X"00040004000004250800E900000604000400000808F4210C1104230F2B000800",
INIT_13 => X"13001A00259000F8F4040400F3000009F8F4040400072B250D90F49000350008",
INIT_14 => X"080401000000000800E600252525000400040004000810210008000E2100080C",
INIT_15 => X"1414242704140100081825040118182427041801000810242710102504011024",
INIT_16 => X"00080002000800000100080C0000081C2504011C1C2427041C01000814250401",
INIT_17 => X"0000006E0068005E0000080C000800240402FB030000080025C007000024C700",
INIT_18 => X"00000008002400000020DF000008002400000010EF0000080024F70000080008",
INIT_19 => X"000905250A1418401008080009071C080400252825982025142E181C240420D8",
INIT_1A => X"980008000A020C14402510259A04054098000C000E01010125030114010C0408",
INIT_1B => X"D400030F257EC4001A00042525741C1418E0280814181C20252410184008F140",
INIT_1C => X"2B211018FF0C000820082514181C20201825141C0200080104257E5C0008257E",
INIT_1D => X"25000225F5001C21019825FF0B000025142525E80008251C0201080010012509",
INIT_1E => X"041021020008010C0008251C020008000C0125042B210C14000C000418080014",
INIT_1F => X"2121001800060008001321140C00180004102100100005000802100026002600",
INIT_20 => X"00100820D825251425181C2509181C140704E00000080C212100140006000410",
INIT_21 => X"2514009A00009A08009A04000707040000250C1410E800F501B300000000F32B",
INIT_22 => X"01F5FFFF01000000082A23232521FF254414E8230801FB000300002500189A10",
INIT_23 => X"0000254D002100022D210525F5FF0312301021010D1A020A252326C318080014",
INIT_24 => X"571014E8006200370008FFFC01FF01252525080108232BFFFF01F80109000500",
INIT_25 => X"08141825081C2550FF14181CE020081418081C25502514181CE0180810081425",
INIT_26 => X"0825500004000D00000D0A252520241014181CD81808FF10140825571410E820",
INIT_27 => X"D40B0600EC0B0200140B181CF025E0000028081014181C202400F1082550FF01",
INIT_28 => X"680000D86ED40000D4680000C86EC4000000014C300B1F00440B0800540B0700",
INIT_29 => X"2020D420070CDC1008D71010D4105F0CDC0008D700D0D400130050001400FED0",
INIT_2A => X"181CA08F000000F88F008400E8AC00D4006800F40101EB0004E0000CDC2008D7",
INIT_2B => X"3030004E20650030702F0000742F000065002020002020004E41564520082514",
INIT_2C => X"000090900000F8A000006F2F00302F00336E2F00326E2F00316E2F00306E2F00",
INIT_2D => X"00744C5245696975652E7468010075000008540000089000000090900000F8A0",
INIT_2E => X"00089000A00002070B000000000000000000000074722E2E4173006474690064",
INIT_2F => X"74722E2E417300647469006400744C5245696975652E74680100750000085400",
INIT_30 => X"2A0001000020200000011E0004000024A00002070B0000000000000000000000",
INIT_31 => X"0301420001000020006003083801040000D030903201300010000060D0300701",
INIT_32 => X"00000000530001000000207003084D00100000D020A003084800100000200080",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic