---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"8E3CAF273C14AC2C008C3C00088C3C24088C3C3C000000000003273C0003273C",
INIT_01 => X"008C3C27038F8F2408AC8C3C3CAE10001428008E000CAC24AF3C8C0024AE243C",
INIT_02 => X"3CAC24ACAC003C2400340003000327083C8F240C3C8C3C3C0C3C0CAF27001030",
INIT_03 => X"243C243C241400AC243C243C241400AC243C243C273C273C000000030014008C",
INIT_04 => X"AFAFAFAFAFAFAFAF2308000C24142400AC8C243C243C243C24142400AC8C243C",
INIT_05 => X"8F230CAF0008200010002000108C3CAF00AF00AF2340AFAFAFAFAFAFAFAFAFAF",
INIT_06 => X"3423038F038F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F0008ACAC3C0020",
INIT_07 => X"0003AC00008CAC34248C0003001030008C0003001030008C0000004003404003",
INIT_08 => X"240024300003AC3C3400033C13008C00243C00240003AC00248C0003AC34008C",
INIT_09 => X"0000000003AC00308CAC00008CAC0030008CAC00008CAC00008C3CAC00243C00",
INIT_0A => X"248C0003AC00248C0003AC34008C0008000800080003AC340003ACAC340003AC",
INIT_0B => X"10240C00AF10AFAF3230AF2700000003AC00008CAC34248C0003AC00008CAC34",
INIT_0C => X"27038F8F8F028FAEAE10240C001232AE0010020CAE14240C001032ACACACAC00",
INIT_0D => X"00250C013010008100AF000027000300AC242403A0AC24001000248C3010008C",
INIT_0E => X"8E92001002008E00AFAF8CAF270003AC240014008C2703008F0000100010008D",
INIT_0F => X"0CAFAF270008000800000027088F028F000CAFAF2727038FAE8F8F8E0010260C",
INIT_10 => X"038F8F00AE8F000C00AFAFAF2727038F8FAE8F000C00AFAFAF2727038F8E8F00",
INIT_11 => X"26AE020C00140010008224240000AFAFAFAFAFAF2727038F8E8F000CAFAF2727",
INIT_12 => X"240C243CAF0CAFAF2424273C00030003000027038F8F8F8F8F8F0010AE020C82",
INIT_13 => X"2724AF3CAF0CAEAF273CAF2627AF3C27AF27AF273C0C240C240C243C240C243C",
INIT_14 => X"3C360C24360C24260C243C360C24360C24260C243C3C0CAF0CAFAFAC3C3CAFAF",
INIT_15 => X"6F4821540A4F4C49004F4C4921544953410010240C8E3C360C24360C24260C34",
INIT_16 => X"547361742E612E65455443646C2E2E6E61730000000F410003273C0000000049",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000075747500",
INIT_18 => X"2E612E65455443646C2E2E6E61730000000F410003273C000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000007574750054736174",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"00000000006F0000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"0310B0BD0440644400620300004402A5004405020000000000405A1A00405A1A",
INIT_01 => X"004202BDE0B0BFA5004084050200000040420002000043A5BF02846202026205",
INIT_02 => X"0343034344000203820200E000E0BD0004BFA50005440204000400BFBD004042",
INIT_03 => X"A505C606A560A4A08404A505A560A4A08404A505BD1D9C1C000000E000400062",
INIT_04 => X"A8A7A6A5A4A3A2A1BD000000A560C6A4A3C38404A505C606A560C6A4A3C38404",
INIT_05 => X"A4A500A400008406A8C5050006C606BB00BB00BA5A1ABFB9B8AFAEADACABAAA9",
INIT_06 => X"1BBD60BB60BBBABFB9B8AFAEADACABAAA9A8A7A6A5A4A3A2A10000C0C5068505",
INIT_07 => X"00E0824300828242038200E0004042008200E0004042008200000084E0029B40",
INIT_08 => X"424303A200E0430263002003200099448404048400E08243038200E082420082",
INIT_09 => X"00000000E045A3A54343640544448684054644830344446400440244C2420202",
INIT_0A => X"038200E08243038200E08242008200000000000000E085A500E08582A200E085",
INIT_0B => X"40040080B040B2BF22B1B1BD000000E0824300828242038200E0824300828242",
INIT_0C => X"BDE0B0B1B200BF02024004000020310200000000024004000040224040405240",
INIT_0D => X"E2080020A5A0000500BFA080BD00E000820202E0C582C20060C24286A5400082",
INIT_0E => X"0425004022000280BFB091B1BD00E0820200400082BDE000BF000000E0400022",
INIT_0F => X"00B0BFBD00000000000000BD00B000BF8000BFB0BDBDE0B002B1BF0200003100",
INIT_10 => X"E0B0B10011BF8000A0B0B1BFBDBDE0B0B111BF8000A0B0B1BFBDBDE0B002BF80",
INIT_11 => X"103320000052004000021312A080B4BFB0B1B2B3BDBDE0B002BF8000B0BFBDBD",
INIT_12 => X"84000504B000B1BF8405BD0400E000E00000BDE0B0B1B2B3B4BF000034200014",
INIT_13 => X"A342A202A00022A4A211A204A2A210A2A2A2A2A2040004008400050484000504",
INIT_14 => X"050400050400050400A5050400050400050400A5050400A000A0A0430204A2A2",
INIT_15 => X"2065006500464552004E45520D494F53430000A50024050400050400050400A5",
INIT_16 => X"4173006469747278004154006462676F62742E0701670000405A1A000000004E",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000074722E2E",
INIT_18 => X"69747278004154006462676F62742E0701670000405A1A000000000000000000",
INIT_19 => X"00000000000000000000000000000000000000000000000074722E2E41730064",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000FF0000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"0B0000FF00000B00000B0000010B000A010B0000000000000000020000000100",
INIT_01 => X"000040000000000A01030B00200B00000000000B0001030A00200B18000B0000",
INIT_02 => X"200200020220200000C300000000000140000A01000B004000400100FF000000",
INIT_03 => X"0B000A0000FF18000B000B0000FF18000C000B000E000B000000000000FF0002",
INIT_04 => X"0000000000000000FF00000200FF001800000B000B000A0000FF001800000B00",
INIT_05 => X"00000100000000300040002000002000D800D800FF7000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000202800",
INIT_07 => X"0000001000000000FF00000000FF000000000000FF0000000000006000606000",
INIT_08 => X"0018000000000320BE0000DE000000200B00100000000010FF00000000000000",
INIT_09 => X"00000000000028000000182C00002000240000201800002000002000100B0030",
INIT_0A => X"FF0000000010FF00000000000000000100010000000000000000000000000000",
INIT_0B => X"0000019000000000000000FF00000000001000000000FF000000001000000000",
INIT_0C => X"000000000010000000FF00010000000080002001000000010000000000000080",
INIT_0D => X"380001200000000038004048FF00001000000000000000100018000000000000",
INIT_0E => X"000000001000008000000000FF10000000000000000000000010000010FF0000",
INIT_0F => X"000000FF00020002000000000100200080010000FF0000000000000000FF0002",
INIT_10 => X"000000100000800088000000FF000000000000800088000000FF000000000080",
INIT_11 => X"0000200000000000000000008088000000000000FF000000000080000000FF00",
INIT_12 => X"00010000000100000000FF00000010000000000000000000000000FF002000FF",
INIT_13 => X"0000004000010B00000000010000200000000000400100000001000000010000",
INIT_14 => X"0002010002010002014B000201000201000201651D4001000100000B00400000",
INIT_15 => X"4D6C007300464443000D44430A4F4C204300FF0A010B000201000201000201A1",
INIT_16 => X"43002E616E616F742E424F562D756E7400727304006E0000000200000000000A",
INIT_17 => X"00000B0000000000000000000000000000000000000000000000000065696167",
INIT_18 => X"6E616F742E424F562D756E7400727304006E0000000200000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000006569616743002E61",
INIT_1A => X"0B0A00000000000000000B0A000000000000000A000000000000000000000B00",
INIT_1B => X"00000B0000FF0000000000020B0C00000000000000010B0B0000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000B00000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"1C0010E80018180100180000D31400BCB31400000000000000085C000008A000",
INIT_01 => X"00040018081014E0B3081400001C07000907001C00B308D014001404011C0100",
INIT_02 => X"00000A000C120009185000080008185E0014F0B300100000E8006814E8001001",
INIT_03 => X"1000C00004FD2A001000100004FD2A0020001000200010000000000800FD0008",
INIT_04 => X"2C2824201C1814109896005404FB042A000010001000BC0004FB042A00001000",
INIT_05 => X"64000C6400B601420424012013080060125C1058FC0054504C4844403C383430",
INIT_06 => X"01681360115C5854504C4844403C3834302C2824201C18141000B21010000401",
INIT_07 => X"0008002400000001FE00000800FC020004000800FC0100040000000008000008",
INIT_08 => X"2004011F00080800EF0008AD030000212000802000080024FD00000800020000",
INIT_09 => X"00000000081C25011C1C24421C14250102141424271418250018000021200080",
INIT_0A => X"EF0000080024F7000008000800000006000000F600080002000800000100080C",
INIT_0B => X"0E18F8251013181C03FF14E000000008002400000020DF000008002400000010",
INIT_0C => X"2008101418251C1008F540F80006020C250A25FA040540F8000A011408040025",
INIT_0D => X"2101A025FF0B000025142525E80008251402010800100125092B4010FF0B0008",
INIT_0E => X"000000072B0010251C140818E025081402000300081808001425000225F50014",
INIT_0F => X"EF1014E80052005000000018FA10251425D31410E820081410181C0800F60113",
INIT_10 => X"08141825081C25E82514181CE020081418081C25E82514181CE0180810081425",
INIT_11 => X"010825E80004000D00000D0A252520241014181CD8180810081425EF1014E820",
INIT_12 => X"541C0300C41CC8CCF402300000082508000028081014181C202400F10825E8FF",
INIT_13 => X"90089000BC0014A8A800B80050B40010B050AC10005E01E2301C1F00441C0400",
INIT_14 => X"0710480C1043081040404C00480C004308004000CD0052A4009C94100000A098",
INIT_15 => X"416C0074000D2020000A2020004E41564500FFF8B3140020480C204308204020",
INIT_16 => X"4B53627469006400744C5245696975652E74680100750000085C000000000000",
INIT_17 => X"0020A40000011E0004000024A00002070B00000000000000000000007362746E",
INIT_18 => X"69006400744C5245696975652E74680100750000085C0000D03007012A000100",
INIT_19 => X"00011E0004000024A00002070B00000000000000000000007362746E4B536274",
INIT_1A => X"C4BC01013801040000485CBC320130001000008CD03007012A0001000020A400",
INIT_1B => X"0010C40000F54D0001000000B0200308470010000010B0100308420001000000",
INIT_1C => X"000000000000000000000000000000000000000000000000D400000301000100",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic