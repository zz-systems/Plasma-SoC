// de1_soc.v

// Generated using ACDS version 13.1 162 at 2018.09.10.21:24:01

`timescale 1 ps / 1 ps
module de1_soc (
		input  wire        clk_clk,                             //                          clk.clk
		output wire [6:0]  hex_0_external_connection_export,    //    hex_0_external_connection.export
		output wire [6:0]  hex_1_external_connection_export,    //    hex_1_external_connection.export
		output wire [6:0]  hex_2_external_connection_export,    //    hex_2_external_connection.export
		output wire [6:0]  hex_3_external_connection_export,    //    hex_3_external_connection.export
		output wire [6:0]  hex_4_external_connection_export,    //    hex_4_external_connection.export
		output wire [6:0]  hex_5_external_connection_export,    //    hex_5_external_connection.export
		output wire [14:0] hps_0_ddr_mem_a,                     //                    hps_0_ddr.mem_a
		output wire [2:0]  hps_0_ddr_mem_ba,                    //                             .mem_ba
		output wire        hps_0_ddr_mem_ck,                    //                             .mem_ck
		output wire        hps_0_ddr_mem_ck_n,                  //                             .mem_ck_n
		output wire        hps_0_ddr_mem_cke,                   //                             .mem_cke
		output wire        hps_0_ddr_mem_cs_n,                  //                             .mem_cs_n
		output wire        hps_0_ddr_mem_ras_n,                 //                             .mem_ras_n
		output wire        hps_0_ddr_mem_cas_n,                 //                             .mem_cas_n
		output wire        hps_0_ddr_mem_we_n,                  //                             .mem_we_n
		output wire        hps_0_ddr_mem_reset_n,               //                             .mem_reset_n
		inout  wire [31:0] hps_0_ddr_mem_dq,                    //                             .mem_dq
		inout  wire [3:0]  hps_0_ddr_mem_dqs,                   //                             .mem_dqs
		inout  wire [3:0]  hps_0_ddr_mem_dqs_n,                 //                             .mem_dqs_n
		output wire        hps_0_ddr_mem_odt,                   //                             .mem_odt
		output wire [3:0]  hps_0_ddr_mem_dm,                    //                             .mem_dm
		input  wire        hps_0_ddr_oct_rzqin,                 //                             .oct_rzqin
		output wire        hps_io_0_hps_io_emac1_inst_TX_CLK,   //                     hps_io_0.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_0_hps_io_emac1_inst_TXD0,     //                             .hps_io_emac1_inst_TXD0
		output wire        hps_io_0_hps_io_emac1_inst_TXD1,     //                             .hps_io_emac1_inst_TXD1
		output wire        hps_io_0_hps_io_emac1_inst_TXD2,     //                             .hps_io_emac1_inst_TXD2
		output wire        hps_io_0_hps_io_emac1_inst_TXD3,     //                             .hps_io_emac1_inst_TXD3
		input  wire        hps_io_0_hps_io_emac1_inst_RXD0,     //                             .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_0_hps_io_emac1_inst_MDIO,     //                             .hps_io_emac1_inst_MDIO
		output wire        hps_io_0_hps_io_emac1_inst_MDC,      //                             .hps_io_emac1_inst_MDC
		input  wire        hps_io_0_hps_io_emac1_inst_RX_CTL,   //                             .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_0_hps_io_emac1_inst_TX_CTL,   //                             .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_0_hps_io_emac1_inst_RX_CLK,   //                             .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_0_hps_io_emac1_inst_RXD1,     //                             .hps_io_emac1_inst_RXD1
		input  wire        hps_io_0_hps_io_emac1_inst_RXD2,     //                             .hps_io_emac1_inst_RXD2
		input  wire        hps_io_0_hps_io_emac1_inst_RXD3,     //                             .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_0_hps_io_qspi_inst_IO0,       //                             .hps_io_qspi_inst_IO0
		inout  wire        hps_io_0_hps_io_qspi_inst_IO1,       //                             .hps_io_qspi_inst_IO1
		inout  wire        hps_io_0_hps_io_qspi_inst_IO2,       //                             .hps_io_qspi_inst_IO2
		inout  wire        hps_io_0_hps_io_qspi_inst_IO3,       //                             .hps_io_qspi_inst_IO3
		output wire        hps_io_0_hps_io_qspi_inst_SS0,       //                             .hps_io_qspi_inst_SS0
		output wire        hps_io_0_hps_io_qspi_inst_CLK,       //                             .hps_io_qspi_inst_CLK
		inout  wire        hps_io_0_hps_io_sdio_inst_CMD,       //                             .hps_io_sdio_inst_CMD
		inout  wire        hps_io_0_hps_io_sdio_inst_D0,        //                             .hps_io_sdio_inst_D0
		inout  wire        hps_io_0_hps_io_sdio_inst_D1,        //                             .hps_io_sdio_inst_D1
		output wire        hps_io_0_hps_io_sdio_inst_CLK,       //                             .hps_io_sdio_inst_CLK
		inout  wire        hps_io_0_hps_io_sdio_inst_D2,        //                             .hps_io_sdio_inst_D2
		inout  wire        hps_io_0_hps_io_sdio_inst_D3,        //                             .hps_io_sdio_inst_D3
		inout  wire        hps_io_0_hps_io_usb1_inst_D0,        //                             .hps_io_usb1_inst_D0
		inout  wire        hps_io_0_hps_io_usb1_inst_D1,        //                             .hps_io_usb1_inst_D1
		inout  wire        hps_io_0_hps_io_usb1_inst_D2,        //                             .hps_io_usb1_inst_D2
		inout  wire        hps_io_0_hps_io_usb1_inst_D3,        //                             .hps_io_usb1_inst_D3
		inout  wire        hps_io_0_hps_io_usb1_inst_D4,        //                             .hps_io_usb1_inst_D4
		inout  wire        hps_io_0_hps_io_usb1_inst_D5,        //                             .hps_io_usb1_inst_D5
		inout  wire        hps_io_0_hps_io_usb1_inst_D6,        //                             .hps_io_usb1_inst_D6
		inout  wire        hps_io_0_hps_io_usb1_inst_D7,        //                             .hps_io_usb1_inst_D7
		input  wire        hps_io_0_hps_io_usb1_inst_CLK,       //                             .hps_io_usb1_inst_CLK
		output wire        hps_io_0_hps_io_usb1_inst_STP,       //                             .hps_io_usb1_inst_STP
		input  wire        hps_io_0_hps_io_usb1_inst_DIR,       //                             .hps_io_usb1_inst_DIR
		input  wire        hps_io_0_hps_io_usb1_inst_NXT,       //                             .hps_io_usb1_inst_NXT
		output wire        hps_io_0_hps_io_spim1_inst_CLK,      //                             .hps_io_spim1_inst_CLK
		output wire        hps_io_0_hps_io_spim1_inst_MOSI,     //                             .hps_io_spim1_inst_MOSI
		input  wire        hps_io_0_hps_io_spim1_inst_MISO,     //                             .hps_io_spim1_inst_MISO
		output wire        hps_io_0_hps_io_spim1_inst_SS0,      //                             .hps_io_spim1_inst_SS0
		input  wire        hps_io_0_hps_io_uart0_inst_RX,       //                             .hps_io_uart0_inst_RX
		output wire        hps_io_0_hps_io_uart0_inst_TX,       //                             .hps_io_uart0_inst_TX
		inout  wire        hps_io_0_hps_io_i2c0_inst_SDA,       //                             .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_0_hps_io_i2c0_inst_SCL,       //                             .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_0_hps_io_i2c1_inst_SDA,       //                             .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_0_hps_io_i2c1_inst_SCL,       //                             .hps_io_i2c1_inst_SCL
		output wire [9:0]  plasma_soc_0_leds_ld,                //            plasma_soc_0_leds.ld
		output wire        plasma_soc_0_sd_card_spi_cs,         //         plasma_soc_0_sd_card.spi_cs
		input  wire        plasma_soc_0_sd_card_spi_miso,       //                             .spi_miso
		output wire        plasma_soc_0_sd_card_spi_mosi,       //                             .spi_mosi
		output wire        plasma_soc_0_sd_card_spi_sclk,       //                             .spi_sclk
		input  wire [9:0]  plasma_soc_0_switches_sw,            //        plasma_soc_0_switches.sw
		input  wire        plasma_soc_0_uart_uart_rx,           //            plasma_soc_0_uart.uart_rx
		output wire        plasma_soc_0_uart_uart_tx,           //                             .uart_tx
		output wire [12:0] sdram_controller_0_wire_addr,        //      sdram_controller_0_wire.addr
		output wire [1:0]  sdram_controller_0_wire_ba,          //                             .ba
		output wire        sdram_controller_0_wire_cas_n,       //                             .cas_n
		output wire        sdram_controller_0_wire_cke,         //                             .cke
		output wire        sdram_controller_0_wire_cs_n,        //                             .cs_n
		inout  wire [15:0] sdram_controller_0_wire_dq,          //                             .dq
		output wire [1:0]  sdram_controller_0_wire_dqm,         //                             .dqm
		output wire        sdram_controller_0_wire_ras_n,       //                             .ras_n
		output wire        sdram_controller_0_wire_we_n,        //                             .we_n
		input  wire [9:0]  switches_external_connection_export, // switches_external_connection.export
		output wire        pll_0_sdram_clk_clk,                 //              pll_0_sdram_clk.clk
		input  wire        hps_0_f2h_cold_reset_req_reset_n,    //     hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,   //    hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_warm_reset_req_reset_n,    //     hps_0_f2h_warm_reset_req.reset_n
		input  wire [3:0]  buttons_external_connection_export,  //  buttons_external_connection.export
		input  wire        reset_reset_n,                       //                        reset.reset_n
		output wire        hps_0_h2f_reset_reset_n              //              hps_0_h2f_reset.reset_n
	);

	wire          pll_0_outclk0_clk;                                         // pll_0:outclk_0 -> [buttons:clk, hex_0:clk, hex_1:clk, hex_2:clk, hex_3:clk, hex_4:clk, hex_5:clk, hps_0:f2h_axi_clk, hps_0:h2f_axi_clk, hps_0:h2f_lw_axi_clk, hps_master:clk_clk, mm_interconnect_0:pll_0_outclk0_clk, mm_interconnect_1:pll_0_outclk0_clk, mm_interconnect_2:pll_0_outclk0_clk, mm_interconnect_3:pll_0_outclk0_clk, plasma_master:clk_clk, plasma_soc_0:GCLK, rst_controller:clk, rst_controller_002:clk, sdram_controller_0:clk, switches:clk, sysid_qsys_0:clock]
	wire          mm_interconnect_0_sdram_controller_0_s1_waitrequest;       // sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	wire   [15:0] mm_interconnect_0_sdram_controller_0_s1_writedata;         // mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	wire   [24:0] mm_interconnect_0_sdram_controller_0_s1_address;           // mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	wire          mm_interconnect_0_sdram_controller_0_s1_chipselect;        // mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	wire          mm_interconnect_0_sdram_controller_0_s1_write;             // mm_interconnect_0:sdram_controller_0_s1_write -> sdram_controller_0:az_wr_n
	wire          mm_interconnect_0_sdram_controller_0_s1_read;              // mm_interconnect_0:sdram_controller_0_s1_read -> sdram_controller_0:az_rd_n
	wire   [15:0] mm_interconnect_0_sdram_controller_0_s1_readdata;          // sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	wire          mm_interconnect_0_sdram_controller_0_s1_readdatavalid;     // sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	wire    [1:0] mm_interconnect_0_sdram_controller_0_s1_byteenable;        // mm_interconnect_0:sdram_controller_0_s1_byteenable -> sdram_controller_0:az_be_n
	wire    [1:0] plasma_soc_0_avalon_master_0_response;                     // mm_interconnect_0:plasma_soc_0_avalon_master_0_response -> plasma_soc_0:avm_response
	wire          plasma_soc_0_avalon_master_0_waitrequest;                  // mm_interconnect_0:plasma_soc_0_avalon_master_0_waitrequest -> plasma_soc_0:avm_waitrequest_n
	wire   [31:0] plasma_soc_0_avalon_master_0_writedata;                    // plasma_soc_0:avm_writedata -> mm_interconnect_0:plasma_soc_0_avalon_master_0_writedata
	wire   [31:0] plasma_soc_0_avalon_master_0_address;                      // plasma_soc_0:avm_address -> mm_interconnect_0:plasma_soc_0_avalon_master_0_address
	wire          plasma_soc_0_avalon_master_0_write;                        // plasma_soc_0:avm_write -> mm_interconnect_0:plasma_soc_0_avalon_master_0_write
	wire          plasma_soc_0_avalon_master_0_read;                         // plasma_soc_0:avm_read -> mm_interconnect_0:plasma_soc_0_avalon_master_0_read
	wire   [31:0] plasma_soc_0_avalon_master_0_readdata;                     // mm_interconnect_0:plasma_soc_0_avalon_master_0_readdata -> plasma_soc_0:avm_readdata
	wire    [3:0] plasma_soc_0_avalon_master_0_byteenable;                   // plasma_soc_0:avm_byteenable -> mm_interconnect_0:plasma_soc_0_avalon_master_0_byteenable
	wire   [31:0] mm_interconnect_0_hex_0_s1_writedata;                      // mm_interconnect_0:hex_0_s1_writedata -> hex_0:writedata
	wire    [1:0] mm_interconnect_0_hex_0_s1_address;                        // mm_interconnect_0:hex_0_s1_address -> hex_0:address
	wire          mm_interconnect_0_hex_0_s1_chipselect;                     // mm_interconnect_0:hex_0_s1_chipselect -> hex_0:chipselect
	wire          mm_interconnect_0_hex_0_s1_write;                          // mm_interconnect_0:hex_0_s1_write -> hex_0:write_n
	wire   [31:0] mm_interconnect_0_hex_0_s1_readdata;                       // hex_0:readdata -> mm_interconnect_0:hex_0_s1_readdata
	wire   [31:0] mm_interconnect_0_hex_1_s1_writedata;                      // mm_interconnect_0:hex_1_s1_writedata -> hex_1:writedata
	wire    [1:0] mm_interconnect_0_hex_1_s1_address;                        // mm_interconnect_0:hex_1_s1_address -> hex_1:address
	wire          mm_interconnect_0_hex_1_s1_chipselect;                     // mm_interconnect_0:hex_1_s1_chipselect -> hex_1:chipselect
	wire          mm_interconnect_0_hex_1_s1_write;                          // mm_interconnect_0:hex_1_s1_write -> hex_1:write_n
	wire   [31:0] mm_interconnect_0_hex_1_s1_readdata;                       // hex_1:readdata -> mm_interconnect_0:hex_1_s1_readdata
	wire   [31:0] mm_interconnect_0_hex_4_s1_writedata;                      // mm_interconnect_0:hex_4_s1_writedata -> hex_4:writedata
	wire    [1:0] mm_interconnect_0_hex_4_s1_address;                        // mm_interconnect_0:hex_4_s1_address -> hex_4:address
	wire          mm_interconnect_0_hex_4_s1_chipselect;                     // mm_interconnect_0:hex_4_s1_chipselect -> hex_4:chipselect
	wire          mm_interconnect_0_hex_4_s1_write;                          // mm_interconnect_0:hex_4_s1_write -> hex_4:write_n
	wire   [31:0] mm_interconnect_0_hex_4_s1_readdata;                       // hex_4:readdata -> mm_interconnect_0:hex_4_s1_readdata
	wire   [31:0] mm_interconnect_0_buttons_s1_writedata;                    // mm_interconnect_0:buttons_s1_writedata -> buttons:writedata
	wire    [1:0] mm_interconnect_0_buttons_s1_address;                      // mm_interconnect_0:buttons_s1_address -> buttons:address
	wire          mm_interconnect_0_buttons_s1_chipselect;                   // mm_interconnect_0:buttons_s1_chipselect -> buttons:chipselect
	wire          mm_interconnect_0_buttons_s1_write;                        // mm_interconnect_0:buttons_s1_write -> buttons:write_n
	wire   [31:0] mm_interconnect_0_buttons_s1_readdata;                     // buttons:readdata -> mm_interconnect_0:buttons_s1_readdata
	wire   [31:0] mm_interconnect_0_hex_3_s1_writedata;                      // mm_interconnect_0:hex_3_s1_writedata -> hex_3:writedata
	wire    [1:0] mm_interconnect_0_hex_3_s1_address;                        // mm_interconnect_0:hex_3_s1_address -> hex_3:address
	wire          mm_interconnect_0_hex_3_s1_chipselect;                     // mm_interconnect_0:hex_3_s1_chipselect -> hex_3:chipselect
	wire          mm_interconnect_0_hex_3_s1_write;                          // mm_interconnect_0:hex_3_s1_write -> hex_3:write_n
	wire   [31:0] mm_interconnect_0_hex_3_s1_readdata;                       // hex_3:readdata -> mm_interconnect_0:hex_3_s1_readdata
	wire   [31:0] mm_interconnect_0_hex_5_s1_writedata;                      // mm_interconnect_0:hex_5_s1_writedata -> hex_5:writedata
	wire    [1:0] mm_interconnect_0_hex_5_s1_address;                        // mm_interconnect_0:hex_5_s1_address -> hex_5:address
	wire          mm_interconnect_0_hex_5_s1_chipselect;                     // mm_interconnect_0:hex_5_s1_chipselect -> hex_5:chipselect
	wire          mm_interconnect_0_hex_5_s1_write;                          // mm_interconnect_0:hex_5_s1_write -> hex_5:write_n
	wire   [31:0] mm_interconnect_0_hex_5_s1_readdata;                       // hex_5:readdata -> mm_interconnect_0:hex_5_s1_readdata
	wire   [31:0] mm_interconnect_0_hex_2_s1_writedata;                      // mm_interconnect_0:hex_2_s1_writedata -> hex_2:writedata
	wire    [1:0] mm_interconnect_0_hex_2_s1_address;                        // mm_interconnect_0:hex_2_s1_address -> hex_2:address
	wire          mm_interconnect_0_hex_2_s1_chipselect;                     // mm_interconnect_0:hex_2_s1_chipselect -> hex_2:chipselect
	wire          mm_interconnect_0_hex_2_s1_write;                          // mm_interconnect_0:hex_2_s1_write -> hex_2:write_n
	wire   [31:0] mm_interconnect_0_hex_2_s1_readdata;                       // hex_2:readdata -> mm_interconnect_0:hex_2_s1_readdata
	wire   [31:0] mm_interconnect_0_switches_s1_writedata;                   // mm_interconnect_0:switches_s1_writedata -> switches:writedata
	wire    [1:0] mm_interconnect_0_switches_s1_address;                     // mm_interconnect_0:switches_s1_address -> switches:address
	wire          mm_interconnect_0_switches_s1_chipselect;                  // mm_interconnect_0:switches_s1_chipselect -> switches:chipselect
	wire          mm_interconnect_0_switches_s1_write;                       // mm_interconnect_0:switches_s1_write -> switches:write_n
	wire   [31:0] mm_interconnect_0_switches_s1_readdata;                    // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire          hps_0_h2f_lw_axi_master_awvalid;                           // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                            // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                            // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                           // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire          hps_0_h2f_lw_axi_master_arready;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                              // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire          hps_0_h2f_lw_axi_master_rready;                            // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire          hps_0_h2f_lw_axi_master_bready;                            // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                            // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                            // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire          hps_0_h2f_lw_axi_master_arvalid;                           // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                            // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                             // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire          hps_0_h2f_lw_axi_master_awready;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                              // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire          hps_0_h2f_lw_axi_master_bvalid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                               // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                            // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                           // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                             // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_rvalid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                             // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_wready;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                           // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                            // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                           // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                             // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                            // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_wvalid;                            // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire          hps_0_h2f_lw_axi_master_wlast;                             // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire          hps_0_h2f_lw_axi_master_rlast;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire    [0:0] mm_interconnect_1_sysid_qsys_0_control_slave_address;      // mm_interconnect_1:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [31:0] mm_interconnect_1_sysid_qsys_0_control_slave_readdata;     // sysid_qsys_0:readdata -> mm_interconnect_1:sysid_qsys_0_control_slave_readdata
	wire          plasma_master_master_waitrequest;                          // mm_interconnect_2:plasma_master_master_waitrequest -> plasma_master:master_waitrequest
	wire   [31:0] plasma_master_master_writedata;                            // plasma_master:master_writedata -> mm_interconnect_2:plasma_master_master_writedata
	wire   [31:0] plasma_master_master_address;                              // plasma_master:master_address -> mm_interconnect_2:plasma_master_master_address
	wire          plasma_master_master_write;                                // plasma_master:master_write -> mm_interconnect_2:plasma_master_master_write
	wire          plasma_master_master_read;                                 // plasma_master:master_read -> mm_interconnect_2:plasma_master_master_read
	wire   [31:0] plasma_master_master_readdata;                             // mm_interconnect_2:plasma_master_master_readdata -> plasma_master:master_readdata
	wire    [3:0] plasma_master_master_byteenable;                           // plasma_master:master_byteenable -> mm_interconnect_2:plasma_master_master_byteenable
	wire          plasma_master_master_readdatavalid;                        // mm_interconnect_2:plasma_master_master_readdatavalid -> plasma_master:master_readdatavalid
	wire          hps_0_h2f_axi_master_awvalid;                              // hps_0:h2f_AWVALID -> mm_interconnect_2:hps_0_h2f_axi_master_awvalid
	wire    [2:0] hps_0_h2f_axi_master_arsize;                               // hps_0:h2f_ARSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_arsize
	wire    [1:0] hps_0_h2f_axi_master_arlock;                               // hps_0:h2f_ARLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_arlock
	wire    [3:0] hps_0_h2f_axi_master_awcache;                              // hps_0:h2f_AWCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_awcache
	wire          hps_0_h2f_axi_master_arready;                              // mm_interconnect_2:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [11:0] hps_0_h2f_axi_master_arid;                                 // hps_0:h2f_ARID -> mm_interconnect_2:hps_0_h2f_axi_master_arid
	wire          hps_0_h2f_axi_master_rready;                               // hps_0:h2f_RREADY -> mm_interconnect_2:hps_0_h2f_axi_master_rready
	wire          hps_0_h2f_axi_master_bready;                               // hps_0:h2f_BREADY -> mm_interconnect_2:hps_0_h2f_axi_master_bready
	wire    [2:0] hps_0_h2f_axi_master_awsize;                               // hps_0:h2f_AWSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_awsize
	wire    [2:0] hps_0_h2f_axi_master_awprot;                               // hps_0:h2f_AWPROT -> mm_interconnect_2:hps_0_h2f_axi_master_awprot
	wire          hps_0_h2f_axi_master_arvalid;                              // hps_0:h2f_ARVALID -> mm_interconnect_2:hps_0_h2f_axi_master_arvalid
	wire    [2:0] hps_0_h2f_axi_master_arprot;                               // hps_0:h2f_ARPROT -> mm_interconnect_2:hps_0_h2f_axi_master_arprot
	wire   [11:0] hps_0_h2f_axi_master_bid;                                  // mm_interconnect_2:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                // hps_0:h2f_ARLEN -> mm_interconnect_2:hps_0_h2f_axi_master_arlen
	wire          hps_0_h2f_axi_master_awready;                              // mm_interconnect_2:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [11:0] hps_0_h2f_axi_master_awid;                                 // hps_0:h2f_AWID -> mm_interconnect_2:hps_0_h2f_axi_master_awid
	wire          hps_0_h2f_axi_master_bvalid;                               // mm_interconnect_2:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [11:0] hps_0_h2f_axi_master_wid;                                  // hps_0:h2f_WID -> mm_interconnect_2:hps_0_h2f_axi_master_wid
	wire    [1:0] hps_0_h2f_axi_master_awlock;                               // hps_0:h2f_AWLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_awlock
	wire    [1:0] hps_0_h2f_axi_master_awburst;                              // hps_0:h2f_AWBURST -> mm_interconnect_2:hps_0_h2f_axi_master_awburst
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                // mm_interconnect_2:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                                // hps_0:h2f_WSTRB -> mm_interconnect_2:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_rvalid;                               // mm_interconnect_2:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire  [127:0] hps_0_h2f_axi_master_wdata;                                // hps_0:h2f_WDATA -> mm_interconnect_2:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_wready;                               // mm_interconnect_2:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                              // hps_0:h2f_ARBURST -> mm_interconnect_2:hps_0_h2f_axi_master_arburst
	wire  [127:0] hps_0_h2f_axi_master_rdata;                                // mm_interconnect_2:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire   [29:0] hps_0_h2f_axi_master_araddr;                               // hps_0:h2f_ARADDR -> mm_interconnect_2:hps_0_h2f_axi_master_araddr
	wire    [3:0] hps_0_h2f_axi_master_arcache;                              // hps_0:h2f_ARCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_arcache
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                // hps_0:h2f_AWLEN -> mm_interconnect_2:hps_0_h2f_axi_master_awlen
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                               // hps_0:h2f_AWADDR -> mm_interconnect_2:hps_0_h2f_axi_master_awaddr
	wire   [11:0] hps_0_h2f_axi_master_rid;                                  // mm_interconnect_2:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_wvalid;                               // hps_0:h2f_WVALID -> mm_interconnect_2:hps_0_h2f_axi_master_wvalid
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                // mm_interconnect_2:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire          hps_0_h2f_axi_master_wlast;                                // hps_0:h2f_WLAST -> mm_interconnect_2:hps_0_h2f_axi_master_wlast
	wire          hps_0_h2f_axi_master_rlast;                                // mm_interconnect_2:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire    [1:0] mm_interconnect_2_plasma_soc_0_avalon_slave_0_response;    // plasma_soc_0:avs_response -> mm_interconnect_2:plasma_soc_0_avalon_slave_0_response
	wire          mm_interconnect_2_plasma_soc_0_avalon_slave_0_waitrequest; // plasma_soc_0:avs_waitrequest_n -> mm_interconnect_2:plasma_soc_0_avalon_slave_0_waitrequest
	wire   [31:0] mm_interconnect_2_plasma_soc_0_avalon_slave_0_writedata;   // mm_interconnect_2:plasma_soc_0_avalon_slave_0_writedata -> plasma_soc_0:avs_writedata
	wire   [31:0] mm_interconnect_2_plasma_soc_0_avalon_slave_0_address;     // mm_interconnect_2:plasma_soc_0_avalon_slave_0_address -> plasma_soc_0:avs_address
	wire          mm_interconnect_2_plasma_soc_0_avalon_slave_0_write;       // mm_interconnect_2:plasma_soc_0_avalon_slave_0_write -> plasma_soc_0:avs_write
	wire          mm_interconnect_2_plasma_soc_0_avalon_slave_0_read;        // mm_interconnect_2:plasma_soc_0_avalon_slave_0_read -> plasma_soc_0:avs_read
	wire   [31:0] mm_interconnect_2_plasma_soc_0_avalon_slave_0_readdata;    // plasma_soc_0:avs_readdata -> mm_interconnect_2:plasma_soc_0_avalon_slave_0_readdata
	wire    [3:0] mm_interconnect_2_plasma_soc_0_avalon_slave_0_byteenable;  // mm_interconnect_2:plasma_soc_0_avalon_slave_0_byteenable -> plasma_soc_0:avs_byteenable
	wire          hps_master_master_waitrequest;                             // mm_interconnect_3:hps_master_master_waitrequest -> hps_master:master_waitrequest
	wire   [31:0] hps_master_master_writedata;                               // hps_master:master_writedata -> mm_interconnect_3:hps_master_master_writedata
	wire   [31:0] hps_master_master_address;                                 // hps_master:master_address -> mm_interconnect_3:hps_master_master_address
	wire          hps_master_master_write;                                   // hps_master:master_write -> mm_interconnect_3:hps_master_master_write
	wire          hps_master_master_read;                                    // hps_master:master_read -> mm_interconnect_3:hps_master_master_read
	wire   [31:0] hps_master_master_readdata;                                // mm_interconnect_3:hps_master_master_readdata -> hps_master:master_readdata
	wire    [3:0] hps_master_master_byteenable;                              // hps_master:master_byteenable -> mm_interconnect_3:hps_master_master_byteenable
	wire          hps_master_master_readdatavalid;                           // mm_interconnect_3:hps_master_master_readdatavalid -> hps_master:master_readdatavalid
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_awvalid;             // mm_interconnect_3:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [2:0] mm_interconnect_3_hps_0_f2h_axi_slave_arsize;              // mm_interconnect_3:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire    [1:0] mm_interconnect_3_hps_0_f2h_axi_slave_arlock;              // mm_interconnect_3:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [3:0] mm_interconnect_3_hps_0_f2h_axi_slave_awcache;             // mm_interconnect_3:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_arready;             // hps_0:f2h_ARREADY -> mm_interconnect_3:hps_0_f2h_axi_slave_arready
	wire    [7:0] mm_interconnect_3_hps_0_f2h_axi_slave_arid;                // mm_interconnect_3:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_rready;              // mm_interconnect_3:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_bready;              // mm_interconnect_3:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire    [2:0] mm_interconnect_3_hps_0_f2h_axi_slave_awsize;              // mm_interconnect_3:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire    [2:0] mm_interconnect_3_hps_0_f2h_axi_slave_awprot;              // mm_interconnect_3:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_arvalid;             // mm_interconnect_3:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [2:0] mm_interconnect_3_hps_0_f2h_axi_slave_arprot;              // mm_interconnect_3:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [7:0] mm_interconnect_3_hps_0_f2h_axi_slave_bid;                 // hps_0:f2h_BID -> mm_interconnect_3:hps_0_f2h_axi_slave_bid
	wire    [3:0] mm_interconnect_3_hps_0_f2h_axi_slave_arlen;               // mm_interconnect_3:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_awready;             // hps_0:f2h_AWREADY -> mm_interconnect_3:hps_0_f2h_axi_slave_awready
	wire    [7:0] mm_interconnect_3_hps_0_f2h_axi_slave_awid;                // mm_interconnect_3:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_bvalid;              // hps_0:f2h_BVALID -> mm_interconnect_3:hps_0_f2h_axi_slave_bvalid
	wire    [7:0] mm_interconnect_3_hps_0_f2h_axi_slave_wid;                 // mm_interconnect_3:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [1:0] mm_interconnect_3_hps_0_f2h_axi_slave_awlock;              // mm_interconnect_3:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire    [1:0] mm_interconnect_3_hps_0_f2h_axi_slave_awburst;             // mm_interconnect_3:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [1:0] mm_interconnect_3_hps_0_f2h_axi_slave_bresp;               // hps_0:f2h_BRESP -> mm_interconnect_3:hps_0_f2h_axi_slave_bresp
	wire    [4:0] mm_interconnect_3_hps_0_f2h_axi_slave_aruser;              // mm_interconnect_3:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire    [4:0] mm_interconnect_3_hps_0_f2h_axi_slave_awuser;              // mm_interconnect_3:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire   [15:0] mm_interconnect_3_hps_0_f2h_axi_slave_wstrb;               // mm_interconnect_3:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_rvalid;              // hps_0:f2h_RVALID -> mm_interconnect_3:hps_0_f2h_axi_slave_rvalid
	wire    [1:0] mm_interconnect_3_hps_0_f2h_axi_slave_arburst;             // mm_interconnect_3:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire  [127:0] mm_interconnect_3_hps_0_f2h_axi_slave_wdata;               // mm_interconnect_3:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_wready;              // hps_0:f2h_WREADY -> mm_interconnect_3:hps_0_f2h_axi_slave_wready
	wire  [127:0] mm_interconnect_3_hps_0_f2h_axi_slave_rdata;               // hps_0:f2h_RDATA -> mm_interconnect_3:hps_0_f2h_axi_slave_rdata
	wire   [31:0] mm_interconnect_3_hps_0_f2h_axi_slave_araddr;              // mm_interconnect_3:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [3:0] mm_interconnect_3_hps_0_f2h_axi_slave_arcache;             // mm_interconnect_3:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire    [3:0] mm_interconnect_3_hps_0_f2h_axi_slave_awlen;               // mm_interconnect_3:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire   [31:0] mm_interconnect_3_hps_0_f2h_axi_slave_awaddr;              // mm_interconnect_3:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [7:0] mm_interconnect_3_hps_0_f2h_axi_slave_rid;                 // hps_0:f2h_RID -> mm_interconnect_3:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_wvalid;              // mm_interconnect_3:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire    [1:0] mm_interconnect_3_hps_0_f2h_axi_slave_rresp;               // hps_0:f2h_RRESP -> mm_interconnect_3:hps_0_f2h_axi_slave_rresp
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_wlast;               // mm_interconnect_3:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire          mm_interconnect_3_hps_0_f2h_axi_slave_rlast;               // hps_0:f2h_RLAST -> mm_interconnect_3:hps_0_f2h_axi_slave_rlast
	wire          irq_mapper_receiver0_irq;                                  // switches:irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                  // buttons:irq -> irq_mapper:receiver1_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                        // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                        // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [buttons:reset_n, hex_0:reset_n, hex_1:reset_n, hex_2:reset_n, hex_3:reset_n, hex_4:reset_n, hex_5:reset_n, mm_interconnect_0:plasma_soc_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:sysid_qsys_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:plasma_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:plasma_soc_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_3:hps_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:hps_master_master_translator_reset_reset_bridge_in_reset_reset, plasma_soc_0:RST, sdram_controller_0:reset_n, switches:reset_n, sysid_qsys_0:reset_n]
	wire          rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> pll_0:rst
	wire          rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]

	de1_soc_hex_0 hex_0 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (hex_0_external_connection_export)       // external_connection.export
	);

	de1_soc_hex_0 hex_1 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (hex_1_external_connection_export)       // external_connection.export
	);

	de1_soc_hex_0 hex_2 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (hex_2_external_connection_export)       // external_connection.export
	);

	de1_soc_hex_0 hex_3 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (hex_3_external_connection_export)       // external_connection.export
	);

	de1_soc_hex_0 hex_4 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (hex_4_external_connection_export)       // external_connection.export
	);

	de1_soc_hex_0 hex_5 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (hex_5_external_connection_export)       // external_connection.export
	);

	de1_soc_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (3)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),              //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),             // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),              //  f2h_warm_reset_req.reset_n
		.mem_a                    (hps_0_ddr_mem_a),                               //              memory.mem_a
		.mem_ba                   (hps_0_ddr_mem_ba),                              //                    .mem_ba
		.mem_ck                   (hps_0_ddr_mem_ck),                              //                    .mem_ck
		.mem_ck_n                 (hps_0_ddr_mem_ck_n),                            //                    .mem_ck_n
		.mem_cke                  (hps_0_ddr_mem_cke),                             //                    .mem_cke
		.mem_cs_n                 (hps_0_ddr_mem_cs_n),                            //                    .mem_cs_n
		.mem_ras_n                (hps_0_ddr_mem_ras_n),                           //                    .mem_ras_n
		.mem_cas_n                (hps_0_ddr_mem_cas_n),                           //                    .mem_cas_n
		.mem_we_n                 (hps_0_ddr_mem_we_n),                            //                    .mem_we_n
		.mem_reset_n              (hps_0_ddr_mem_reset_n),                         //                    .mem_reset_n
		.mem_dq                   (hps_0_ddr_mem_dq),                              //                    .mem_dq
		.mem_dqs                  (hps_0_ddr_mem_dqs),                             //                    .mem_dqs
		.mem_dqs_n                (hps_0_ddr_mem_dqs_n),                           //                    .mem_dqs_n
		.mem_odt                  (hps_0_ddr_mem_odt),                             //                    .mem_odt
		.mem_dm                   (hps_0_ddr_mem_dm),                              //                    .mem_dm
		.oct_rzqin                (hps_0_ddr_oct_rzqin),                           //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_0_hps_io_emac1_inst_TX_CLK),             //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_0_hps_io_emac1_inst_TXD0),               //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_0_hps_io_emac1_inst_TXD1),               //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_0_hps_io_emac1_inst_TXD2),               //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_0_hps_io_emac1_inst_TXD3),               //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_0_hps_io_emac1_inst_RXD0),               //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_0_hps_io_emac1_inst_MDIO),               //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_0_hps_io_emac1_inst_MDC),                //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_0_hps_io_emac1_inst_RX_CTL),             //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_0_hps_io_emac1_inst_TX_CTL),             //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_0_hps_io_emac1_inst_RX_CLK),             //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_0_hps_io_emac1_inst_RXD1),               //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_0_hps_io_emac1_inst_RXD2),               //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_0_hps_io_emac1_inst_RXD3),               //                    .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_0_hps_io_qspi_inst_IO0),                 //                    .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_0_hps_io_qspi_inst_IO1),                 //                    .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_0_hps_io_qspi_inst_IO2),                 //                    .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_0_hps_io_qspi_inst_IO3),                 //                    .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_0_hps_io_qspi_inst_SS0),                 //                    .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_0_hps_io_qspi_inst_CLK),                 //                    .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_0_hps_io_sdio_inst_CMD),                 //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_0_hps_io_sdio_inst_D0),                  //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_0_hps_io_sdio_inst_D1),                  //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_0_hps_io_sdio_inst_CLK),                 //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_0_hps_io_sdio_inst_D2),                  //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_0_hps_io_sdio_inst_D3),                  //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_0_hps_io_usb1_inst_D0),                  //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_0_hps_io_usb1_inst_D1),                  //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_0_hps_io_usb1_inst_D2),                  //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_0_hps_io_usb1_inst_D3),                  //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_0_hps_io_usb1_inst_D4),                  //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_0_hps_io_usb1_inst_D5),                  //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_0_hps_io_usb1_inst_D6),                  //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_0_hps_io_usb1_inst_D7),                  //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_0_hps_io_usb1_inst_CLK),                 //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_0_hps_io_usb1_inst_STP),                 //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_0_hps_io_usb1_inst_DIR),                 //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_0_hps_io_usb1_inst_NXT),                 //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_0_hps_io_spim1_inst_CLK),                //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_0_hps_io_spim1_inst_MOSI),               //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_0_hps_io_spim1_inst_MISO),               //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_0_hps_io_spim1_inst_SS0),                //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_0_hps_io_uart0_inst_RX),                 //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_0_hps_io_uart0_inst_TX),                 //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_0_hps_io_i2c0_inst_SDA),                 //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_0_hps_io_i2c0_inst_SCL),                 //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_0_hps_io_i2c1_inst_SDA),                 //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_0_hps_io_i2c1_inst_SCL),                 //                    .hps_io_i2c1_inst_SCL
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //           h2f_reset.reset_n
		.h2f_axi_clk              (pll_0_outclk0_clk),                             //       h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                     //      h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                   //                    .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                    //                    .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                   //                    .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                  //                    .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                   //                    .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                  //                    .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                   //                    .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                  //                    .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                  //                    .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                      //                    .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                    //                    .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                    //                    .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                    //                    .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                   //                    .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                   //                    .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                      //                    .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                    //                    .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                   //                    .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                   //                    .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                     //                    .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                   //                    .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                    //                    .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                   //                    .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                  //                    .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                   //                    .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                  //                    .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                   //                    .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                  //                    .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                  //                    .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                      //                    .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                    //                    .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                    //                    .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                    //                    .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                   //                    .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                   //                    .rready
		.f2h_axi_clk              (pll_0_outclk0_clk),                             //       f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_3_hps_0_f2h_axi_slave_awid),    //       f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_3_hps_0_f2h_axi_slave_awaddr),  //                    .awaddr
		.f2h_AWLEN                (mm_interconnect_3_hps_0_f2h_axi_slave_awlen),   //                    .awlen
		.f2h_AWSIZE               (mm_interconnect_3_hps_0_f2h_axi_slave_awsize),  //                    .awsize
		.f2h_AWBURST              (mm_interconnect_3_hps_0_f2h_axi_slave_awburst), //                    .awburst
		.f2h_AWLOCK               (mm_interconnect_3_hps_0_f2h_axi_slave_awlock),  //                    .awlock
		.f2h_AWCACHE              (mm_interconnect_3_hps_0_f2h_axi_slave_awcache), //                    .awcache
		.f2h_AWPROT               (mm_interconnect_3_hps_0_f2h_axi_slave_awprot),  //                    .awprot
		.f2h_AWVALID              (mm_interconnect_3_hps_0_f2h_axi_slave_awvalid), //                    .awvalid
		.f2h_AWREADY              (mm_interconnect_3_hps_0_f2h_axi_slave_awready), //                    .awready
		.f2h_AWUSER               (mm_interconnect_3_hps_0_f2h_axi_slave_awuser),  //                    .awuser
		.f2h_WID                  (mm_interconnect_3_hps_0_f2h_axi_slave_wid),     //                    .wid
		.f2h_WDATA                (mm_interconnect_3_hps_0_f2h_axi_slave_wdata),   //                    .wdata
		.f2h_WSTRB                (mm_interconnect_3_hps_0_f2h_axi_slave_wstrb),   //                    .wstrb
		.f2h_WLAST                (mm_interconnect_3_hps_0_f2h_axi_slave_wlast),   //                    .wlast
		.f2h_WVALID               (mm_interconnect_3_hps_0_f2h_axi_slave_wvalid),  //                    .wvalid
		.f2h_WREADY               (mm_interconnect_3_hps_0_f2h_axi_slave_wready),  //                    .wready
		.f2h_BID                  (mm_interconnect_3_hps_0_f2h_axi_slave_bid),     //                    .bid
		.f2h_BRESP                (mm_interconnect_3_hps_0_f2h_axi_slave_bresp),   //                    .bresp
		.f2h_BVALID               (mm_interconnect_3_hps_0_f2h_axi_slave_bvalid),  //                    .bvalid
		.f2h_BREADY               (mm_interconnect_3_hps_0_f2h_axi_slave_bready),  //                    .bready
		.f2h_ARID                 (mm_interconnect_3_hps_0_f2h_axi_slave_arid),    //                    .arid
		.f2h_ARADDR               (mm_interconnect_3_hps_0_f2h_axi_slave_araddr),  //                    .araddr
		.f2h_ARLEN                (mm_interconnect_3_hps_0_f2h_axi_slave_arlen),   //                    .arlen
		.f2h_ARSIZE               (mm_interconnect_3_hps_0_f2h_axi_slave_arsize),  //                    .arsize
		.f2h_ARBURST              (mm_interconnect_3_hps_0_f2h_axi_slave_arburst), //                    .arburst
		.f2h_ARLOCK               (mm_interconnect_3_hps_0_f2h_axi_slave_arlock),  //                    .arlock
		.f2h_ARCACHE              (mm_interconnect_3_hps_0_f2h_axi_slave_arcache), //                    .arcache
		.f2h_ARPROT               (mm_interconnect_3_hps_0_f2h_axi_slave_arprot),  //                    .arprot
		.f2h_ARVALID              (mm_interconnect_3_hps_0_f2h_axi_slave_arvalid), //                    .arvalid
		.f2h_ARREADY              (mm_interconnect_3_hps_0_f2h_axi_slave_arready), //                    .arready
		.f2h_ARUSER               (mm_interconnect_3_hps_0_f2h_axi_slave_aruser),  //                    .aruser
		.f2h_RID                  (mm_interconnect_3_hps_0_f2h_axi_slave_rid),     //                    .rid
		.f2h_RDATA                (mm_interconnect_3_hps_0_f2h_axi_slave_rdata),   //                    .rdata
		.f2h_RRESP                (mm_interconnect_3_hps_0_f2h_axi_slave_rresp),   //                    .rresp
		.f2h_RLAST                (mm_interconnect_3_hps_0_f2h_axi_slave_rlast),   //                    .rlast
		.f2h_RVALID               (mm_interconnect_3_hps_0_f2h_axi_slave_rvalid),  //                    .rvalid
		.f2h_RREADY               (mm_interconnect_3_hps_0_f2h_axi_slave_rready),  //                    .rready
		.h2f_lw_axi_clk           (pll_0_outclk0_clk),                             //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                            //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                             //            f2h_irq1.irq
	);

	de1_soc_buttons buttons (
		.clk        (pll_0_outclk0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_buttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buttons_s1_readdata),   //                    .readdata
		.in_port    (buttons_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                 //                 irq.irq
	);

	plasma_soc_top plasma_soc_0 (
		.RST               (rst_controller_reset_out_reset),                            //      reset_sink.reset
		.GCLK              (pll_0_outclk0_clk),                                         //      clock_sink.clk
		.LD                (plasma_soc_0_leds_ld),                                      //            leds.ld
		.SPI_CS            (plasma_soc_0_sd_card_spi_cs),                               //         sd_card.spi_cs
		.SPI_MISO          (plasma_soc_0_sd_card_spi_miso),                             //                .spi_miso
		.SPI_MOSI          (plasma_soc_0_sd_card_spi_mosi),                             //                .spi_mosi
		.SPI_SCLK          (plasma_soc_0_sd_card_spi_sclk),                             //                .spi_sclk
		.SW                (plasma_soc_0_switches_sw),                                  //        switches.sw
		.UART_RX           (plasma_soc_0_uart_uart_rx),                                 //            uart.uart_rx
		.UART_TX           (plasma_soc_0_uart_uart_tx),                                 //                .uart_tx
		.avs_waitrequest_n (mm_interconnect_2_plasma_soc_0_avalon_slave_0_waitrequest), //  avalon_slave_0.waitrequest_n
		.avs_response      (mm_interconnect_2_plasma_soc_0_avalon_slave_0_response),    //                .response
		.avs_address       (mm_interconnect_2_plasma_soc_0_avalon_slave_0_address),     //                .address
		.avs_byteenable    (mm_interconnect_2_plasma_soc_0_avalon_slave_0_byteenable),  //                .byteenable
		.avs_read          (mm_interconnect_2_plasma_soc_0_avalon_slave_0_read),        //                .read
		.avs_readdata      (mm_interconnect_2_plasma_soc_0_avalon_slave_0_readdata),    //                .readdata
		.avs_write         (mm_interconnect_2_plasma_soc_0_avalon_slave_0_write),       //                .write
		.avs_writedata     (mm_interconnect_2_plasma_soc_0_avalon_slave_0_writedata),   //                .writedata
		.avm_waitrequest_n (~plasma_soc_0_avalon_master_0_waitrequest),                 // avalon_master_0.waitrequest_n
		.avm_response      (plasma_soc_0_avalon_master_0_response),                     //                .response
		.avm_address       (plasma_soc_0_avalon_master_0_address),                      //                .address
		.avm_byteenable    (plasma_soc_0_avalon_master_0_byteenable),                   //                .byteenable
		.avm_read          (plasma_soc_0_avalon_master_0_read),                         //                .read
		.avm_readdata      (plasma_soc_0_avalon_master_0_readdata),                     //                .readdata
		.avm_write         (plasma_soc_0_avalon_master_0_write),                        //                .write
		.avm_writedata     (plasma_soc_0_avalon_master_0_writedata)                     //                .writedata
	);

	de1_soc_sdram_controller_0 sdram_controller_0 (
		.clk            (pll_0_outclk0_clk),                                     //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_0_wire_we_n)                           //      .export
	);

	de1_soc_switches switches (
		.clk        (pll_0_outclk0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_switches_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_switches_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_switches_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_switches_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_switches_s1_readdata),   //                    .readdata
		.in_port    (switches_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver0_irq)                  //                 irq.irq
	);

	de1_soc_pll_0 pll_0 (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),                  // outclk0.clk
		.outclk_1 (pll_0_sdram_clk_clk),                // outclk1.clk
		.locked   ()                                    // (terminated)
	);

	de1_soc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_0_outclk0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_0_control_slave_address)   //              .address
	);

	de1_soc_hps_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) hps_master (
		.clk_clk              (pll_0_outclk0_clk),               //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                  //    clk_reset.reset
		.master_address       (hps_master_master_address),       //       master.address
		.master_readdata      (hps_master_master_readdata),      //             .readdata
		.master_read          (hps_master_master_read),          //             .read
		.master_write         (hps_master_master_write),         //             .write
		.master_writedata     (hps_master_master_writedata),     //             .writedata
		.master_waitrequest   (hps_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (hps_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (hps_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                 // master_reset.reset
	);

	de1_soc_hps_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) plasma_master (
		.clk_clk              (pll_0_outclk0_clk),                  //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                     //    clk_reset.reset
		.master_address       (plasma_master_master_address),       //       master.address
		.master_readdata      (plasma_master_master_readdata),      //             .readdata
		.master_read          (plasma_master_master_read),          //             .read
		.master_write         (plasma_master_master_write),         //             .write
		.master_writedata     (plasma_master_master_writedata),     //             .writedata
		.master_waitrequest   (plasma_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (plasma_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (plasma_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                    // master_reset.reset
	);

	de1_soc_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                                   (pll_0_outclk0_clk),                                     //                                 pll_0_outclk0.clk
		.plasma_soc_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // plasma_soc_0_reset_sink_reset_bridge_in_reset.reset
		.plasma_soc_0_avalon_master_0_address                (plasma_soc_0_avalon_master_0_address),                  //                  plasma_soc_0_avalon_master_0.address
		.plasma_soc_0_avalon_master_0_waitrequest            (plasma_soc_0_avalon_master_0_waitrequest),              //                                              .waitrequest
		.plasma_soc_0_avalon_master_0_byteenable             (plasma_soc_0_avalon_master_0_byteenable),               //                                              .byteenable
		.plasma_soc_0_avalon_master_0_read                   (plasma_soc_0_avalon_master_0_read),                     //                                              .read
		.plasma_soc_0_avalon_master_0_readdata               (plasma_soc_0_avalon_master_0_readdata),                 //                                              .readdata
		.plasma_soc_0_avalon_master_0_write                  (plasma_soc_0_avalon_master_0_write),                    //                                              .write
		.plasma_soc_0_avalon_master_0_writedata              (plasma_soc_0_avalon_master_0_writedata),                //                                              .writedata
		.plasma_soc_0_avalon_master_0_response               (plasma_soc_0_avalon_master_0_response),                 //                                              .response
		.buttons_s1_address                                  (mm_interconnect_0_buttons_s1_address),                  //                                    buttons_s1.address
		.buttons_s1_write                                    (mm_interconnect_0_buttons_s1_write),                    //                                              .write
		.buttons_s1_readdata                                 (mm_interconnect_0_buttons_s1_readdata),                 //                                              .readdata
		.buttons_s1_writedata                                (mm_interconnect_0_buttons_s1_writedata),                //                                              .writedata
		.buttons_s1_chipselect                               (mm_interconnect_0_buttons_s1_chipselect),               //                                              .chipselect
		.hex_0_s1_address                                    (mm_interconnect_0_hex_0_s1_address),                    //                                      hex_0_s1.address
		.hex_0_s1_write                                      (mm_interconnect_0_hex_0_s1_write),                      //                                              .write
		.hex_0_s1_readdata                                   (mm_interconnect_0_hex_0_s1_readdata),                   //                                              .readdata
		.hex_0_s1_writedata                                  (mm_interconnect_0_hex_0_s1_writedata),                  //                                              .writedata
		.hex_0_s1_chipselect                                 (mm_interconnect_0_hex_0_s1_chipselect),                 //                                              .chipselect
		.hex_1_s1_address                                    (mm_interconnect_0_hex_1_s1_address),                    //                                      hex_1_s1.address
		.hex_1_s1_write                                      (mm_interconnect_0_hex_1_s1_write),                      //                                              .write
		.hex_1_s1_readdata                                   (mm_interconnect_0_hex_1_s1_readdata),                   //                                              .readdata
		.hex_1_s1_writedata                                  (mm_interconnect_0_hex_1_s1_writedata),                  //                                              .writedata
		.hex_1_s1_chipselect                                 (mm_interconnect_0_hex_1_s1_chipselect),                 //                                              .chipselect
		.hex_2_s1_address                                    (mm_interconnect_0_hex_2_s1_address),                    //                                      hex_2_s1.address
		.hex_2_s1_write                                      (mm_interconnect_0_hex_2_s1_write),                      //                                              .write
		.hex_2_s1_readdata                                   (mm_interconnect_0_hex_2_s1_readdata),                   //                                              .readdata
		.hex_2_s1_writedata                                  (mm_interconnect_0_hex_2_s1_writedata),                  //                                              .writedata
		.hex_2_s1_chipselect                                 (mm_interconnect_0_hex_2_s1_chipselect),                 //                                              .chipselect
		.hex_3_s1_address                                    (mm_interconnect_0_hex_3_s1_address),                    //                                      hex_3_s1.address
		.hex_3_s1_write                                      (mm_interconnect_0_hex_3_s1_write),                      //                                              .write
		.hex_3_s1_readdata                                   (mm_interconnect_0_hex_3_s1_readdata),                   //                                              .readdata
		.hex_3_s1_writedata                                  (mm_interconnect_0_hex_3_s1_writedata),                  //                                              .writedata
		.hex_3_s1_chipselect                                 (mm_interconnect_0_hex_3_s1_chipselect),                 //                                              .chipselect
		.hex_4_s1_address                                    (mm_interconnect_0_hex_4_s1_address),                    //                                      hex_4_s1.address
		.hex_4_s1_write                                      (mm_interconnect_0_hex_4_s1_write),                      //                                              .write
		.hex_4_s1_readdata                                   (mm_interconnect_0_hex_4_s1_readdata),                   //                                              .readdata
		.hex_4_s1_writedata                                  (mm_interconnect_0_hex_4_s1_writedata),                  //                                              .writedata
		.hex_4_s1_chipselect                                 (mm_interconnect_0_hex_4_s1_chipselect),                 //                                              .chipselect
		.hex_5_s1_address                                    (mm_interconnect_0_hex_5_s1_address),                    //                                      hex_5_s1.address
		.hex_5_s1_write                                      (mm_interconnect_0_hex_5_s1_write),                      //                                              .write
		.hex_5_s1_readdata                                   (mm_interconnect_0_hex_5_s1_readdata),                   //                                              .readdata
		.hex_5_s1_writedata                                  (mm_interconnect_0_hex_5_s1_writedata),                  //                                              .writedata
		.hex_5_s1_chipselect                                 (mm_interconnect_0_hex_5_s1_chipselect),                 //                                              .chipselect
		.sdram_controller_0_s1_address                       (mm_interconnect_0_sdram_controller_0_s1_address),       //                         sdram_controller_0_s1.address
		.sdram_controller_0_s1_write                         (mm_interconnect_0_sdram_controller_0_s1_write),         //                                              .write
		.sdram_controller_0_s1_read                          (mm_interconnect_0_sdram_controller_0_s1_read),          //                                              .read
		.sdram_controller_0_s1_readdata                      (mm_interconnect_0_sdram_controller_0_s1_readdata),      //                                              .readdata
		.sdram_controller_0_s1_writedata                     (mm_interconnect_0_sdram_controller_0_s1_writedata),     //                                              .writedata
		.sdram_controller_0_s1_byteenable                    (mm_interconnect_0_sdram_controller_0_s1_byteenable),    //                                              .byteenable
		.sdram_controller_0_s1_readdatavalid                 (mm_interconnect_0_sdram_controller_0_s1_readdatavalid), //                                              .readdatavalid
		.sdram_controller_0_s1_waitrequest                   (mm_interconnect_0_sdram_controller_0_s1_waitrequest),   //                                              .waitrequest
		.sdram_controller_0_s1_chipselect                    (mm_interconnect_0_sdram_controller_0_s1_chipselect),    //                                              .chipselect
		.switches_s1_address                                 (mm_interconnect_0_switches_s1_address),                 //                                   switches_s1.address
		.switches_s1_write                                   (mm_interconnect_0_switches_s1_write),                   //                                              .write
		.switches_s1_readdata                                (mm_interconnect_0_switches_s1_readdata),                //                                              .readdata
		.switches_s1_writedata                               (mm_interconnect_0_switches_s1_writedata),               //                                              .writedata
		.switches_s1_chipselect                              (mm_interconnect_0_switches_s1_chipselect)               //                                              .chipselect
	);

	de1_soc_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                          //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                        //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                         //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                        //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                       //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                        //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                       //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                        //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                       //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                       //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                           //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                         //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                         //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                         //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                        //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                        //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                           //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                         //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                        //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                        //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                          //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                        //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                         //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                        //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                       //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                        //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                       //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                        //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                       //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                       //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                           //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                         //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                         //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                         //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                        //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                        //                                                              .rready
		.pll_0_outclk0_clk                                                   (pll_0_outclk0_clk),                                     //                                                 pll_0_outclk0.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                    // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sysid_qsys_0_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),                        //                      sysid_qsys_0_reset_reset_bridge_in_reset.reset
		.sysid_qsys_0_control_slave_address                                  (mm_interconnect_1_sysid_qsys_0_control_slave_address),  //                                    sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                 (mm_interconnect_1_sysid_qsys_0_control_slave_readdata)  //                                                              .readdata
	);

	de1_soc_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                  //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                 //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                               //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                               //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                               //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                               //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                   //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                 //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                 //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                 //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                   //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                 //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                  //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                 //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                               //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                               //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                               //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                               //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                   //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                 //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                 //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                 //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                //                                                           .rready
		.pll_0_outclk0_clk                                                (pll_0_outclk0_clk),                                          //                                              pll_0_outclk0.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                         // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.plasma_master_clk_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                             //              plasma_master_clk_reset_reset_bridge_in_reset.reset
		.plasma_soc_0_reset_sink_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                             //              plasma_soc_0_reset_sink_reset_bridge_in_reset.reset
		.plasma_master_master_address                                     (plasma_master_master_address),                               //                                       plasma_master_master.address
		.plasma_master_master_waitrequest                                 (plasma_master_master_waitrequest),                           //                                                           .waitrequest
		.plasma_master_master_byteenable                                  (plasma_master_master_byteenable),                            //                                                           .byteenable
		.plasma_master_master_read                                        (plasma_master_master_read),                                  //                                                           .read
		.plasma_master_master_readdata                                    (plasma_master_master_readdata),                              //                                                           .readdata
		.plasma_master_master_readdatavalid                               (plasma_master_master_readdatavalid),                         //                                                           .readdatavalid
		.plasma_master_master_write                                       (plasma_master_master_write),                                 //                                                           .write
		.plasma_master_master_writedata                                   (plasma_master_master_writedata),                             //                                                           .writedata
		.plasma_soc_0_avalon_slave_0_address                              (mm_interconnect_2_plasma_soc_0_avalon_slave_0_address),      //                                plasma_soc_0_avalon_slave_0.address
		.plasma_soc_0_avalon_slave_0_write                                (mm_interconnect_2_plasma_soc_0_avalon_slave_0_write),        //                                                           .write
		.plasma_soc_0_avalon_slave_0_read                                 (mm_interconnect_2_plasma_soc_0_avalon_slave_0_read),         //                                                           .read
		.plasma_soc_0_avalon_slave_0_readdata                             (mm_interconnect_2_plasma_soc_0_avalon_slave_0_readdata),     //                                                           .readdata
		.plasma_soc_0_avalon_slave_0_writedata                            (mm_interconnect_2_plasma_soc_0_avalon_slave_0_writedata),    //                                                           .writedata
		.plasma_soc_0_avalon_slave_0_byteenable                           (mm_interconnect_2_plasma_soc_0_avalon_slave_0_byteenable),   //                                                           .byteenable
		.plasma_soc_0_avalon_slave_0_waitrequest                          (~mm_interconnect_2_plasma_soc_0_avalon_slave_0_waitrequest), //                                                           .waitrequest
		.plasma_soc_0_avalon_slave_0_response                             (mm_interconnect_2_plasma_soc_0_avalon_slave_0_response)      //                                                           .response
	);

	de1_soc_mm_interconnect_3 mm_interconnect_3 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_3_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_3_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_3_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_3_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_3_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_3_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_3_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_3_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_3_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_3_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_3_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_3_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_3_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_3_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_3_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_3_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_3_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_3_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_3_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_3_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_3_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_3_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_3_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_3_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_3_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_3_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_3_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_3_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_3_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_3_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_3_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_3_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_3_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_3_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_3_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_3_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_3_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_3_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.pll_0_outclk0_clk                                                (pll_0_outclk0_clk),                             //                                              pll_0_outclk0.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.hps_master_clk_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                //                 hps_master_clk_reset_reset_bridge_in_reset.reset
		.hps_master_master_translator_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                //   hps_master_master_translator_reset_reset_bridge_in_reset.reset
		.hps_master_master_address                                        (hps_master_master_address),                     //                                          hps_master_master.address
		.hps_master_master_waitrequest                                    (hps_master_master_waitrequest),                 //                                                           .waitrequest
		.hps_master_master_byteenable                                     (hps_master_master_byteenable),                  //                                                           .byteenable
		.hps_master_master_read                                           (hps_master_master_read),                        //                                                           .read
		.hps_master_master_readdata                                       (hps_master_master_readdata),                    //                                                           .readdata
		.hps_master_master_readdatavalid                                  (hps_master_master_readdatavalid),               //                                                           .readdatavalid
		.hps_master_master_write                                          (hps_master_master_write),                       //                                                           .write
		.hps_master_master_writedata                                      (hps_master_master_writedata)                    //                                                           .writedata
	);

	de1_soc_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	de1_soc_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
