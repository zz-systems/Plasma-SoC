---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "text.exe".
--    Run convert.exe to change "text.exe" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "run_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    corectly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"AF27AF24AFAF00001424AC24278C3C24088C3C3C000000000003273C0003273C",
INIT_01 => X"A00093A000932410A0009300108E3C2A020C0000001600000000001400000000",
INIT_02 => X"8E24108EA000938E00102A020C27A00093A000932410A0009300108E2A270C02",
INIT_03 => X"243CAF248E3CAF273C14AC2C008C3C00088C3C27038F8F8F8FA000838EA00083",
INIT_04 => X"243C8E8C3CAF3C2727038F8F8F240824AC3C3CAE1000162A0C24AC24AFAE3C00",
INIT_05 => X"24AC243C1002008E00162402122400300C008C3C001402263CAF14AFAFAFAF00",
INIT_06 => X"3C240CAF3C8E3CAF27001030008C3C27038F8F8F8F8F8FA0AE241200008EA010",
INIT_07 => X"0000000327083C8F8F000C8E240C3C8E240C008E240C3C8E240C008E000C8C8E",
INIT_08 => X"24142400AC8C243C243C243C241400AC243C243C241400AC243C243C273C273C",
INIT_09 => X"AFAFAFAFAFAFAFAFAFAFAFAFAFAF2308000C000C24142400AC8C243C243C243C",
INIT_0A => X"8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F000CAF00AF00AF2340AFAFAFAF",
INIT_0B => X"008CAC34248C0003001030008C0003001030008C0040034040033423038F038F",
INIT_0C => X"14020C24ACAC3C0010240CAFAF00AF270003AC00248C0003AC34008C0003AC00",
INIT_0D => X"2424103C3C14020C2424103C3C14020C24AE1024AE243C3C14020C2424103C3C",
INIT_0E => X"14020C242410AE243C3C14020C242410AE243C3C14020C242410AE3C3C14020C",
INIT_0F => X"AFAFAFAFAF3CAF2700000010000CAF2700000027038F8F028F00020C2410AE3C",
INIT_10 => X"8F8F8F2616263C0C0202000010008E00120014020210028E24243C000026AFAF",
INIT_11 => X"8F028F8F003C0C3002003C0C02AC0024AFAF00240030AF3C2727038F8F8F8F8F",
INIT_12 => X"00008C0010248C3C0024240010AC03ACACAC24AC3C00343C0024243C27083C30",
INIT_13 => X"3C100003ACACACAC008C8C000300108CAC10ACACAC008CACAC240024142C0014",
INIT_14 => X"00008C241000108C008CACACACAC8C00108CAC10ACACAC8C001100001024248C",
INIT_15 => X"00248C000300248C0000000300108C000000ACACACAC008C8CAC2400008C0014",
INIT_16 => X"AC0000308CAC0000008C240003AC0000308CAC0000008C240003AC00008CAC00",
INIT_17 => X"AC00248C0003AC340003ACAC340003AC000003AC0000308CAC0000008C240003",
INIT_18 => X"0003AC34008C000800080008000003AC0003AC00341024108C0003AC0000308C",
INIT_19 => X"AF8CAF2700000003AC00008CAC34248C0003AC00008CAC34248C0003AC00248C",
INIT_1A => X"24AEAE243C16240010AEAE24AEAE243C1624ACACACAC0010000C2400AF12AFAF",
INIT_1B => X"24AE10240C0012001232AEAE240010020CAE14240C00100010322424001024AE",
INIT_1C => X"3C10020C243C2410020C243C10008C00000CAFAFAF2727038F8F8F8F028FAEAE",
INIT_1D => X"AC24001000008C8C3010008C2703008F8F8F27088F028F8F2400102410020C24",
INIT_1E => X"2703008F0000100010008D00250C013010008100AF000027000300AC242403A0",
INIT_1F => X"100014008CAC0010008C2414000300AC24000390AC24001000008C8C0010008C",
INIT_20 => X"10008CAC0000008C0010008C001400108C0010008CAC00008C0010008C241400",
INIT_21 => X"8E001002008E8C270800008F028F8F0014AFAFAF248C278C0003AC0000008C00",
INIT_22 => X"0027088F028F000C8E000C8E000C8E0010248C008E000CAFAF270010260C8C92",
INIT_23 => X"2703008FA01024A02480800010000000000024000CAF27000324100010008000",
INIT_24 => X"1000140080800008A000A1242400040010A11000240000240000152400000000",
INIT_25 => X"8F8E8F000CAFAF27000800080003A01424802400000003340300003030241024",
INIT_26 => X"AFAF2727038F8F00AE8F000C30AFAFAF2727038F8FAE8F000C00AFAFAF272703",
INIT_27 => X"020C9226AE020C00140010008224240000AFAFAFAFAFAF272703308F8F8E000C",
INIT_28 => X"240C243C240C243C240C243CAF0CAFAF2400273C0027038F8F8F8F8F8F0010AE",
INIT_29 => X"0C3C0CAC0C3C3C240C243C3CAE0C263C240C243C3C3C240C240C243C240C243C",
INIT_2A => X"0C36240C36340C263C240C36240C36240C263C240C36240C36240C263C3C0C3C",
INIT_2B => X"2703008F8F8F240C243C3C240C3C8C3C240C3C8E360C360C24240C36240C2624",
INIT_2C => X"7463640030300D4D6C0D006C646477307564723A544F4C494F4C492154495341",
INIT_2D => X"0000000000000000000000007230676400696400746364007463640074636400",
INIT_2E => X"742E612E65455443646C2E2E6E61730000000F410003273C0003273C00000000",
INIT_2F => X"0003273C0003273C0000000000000000000000000000006569616743002E6161",
INIT_30 => X"0000006569616743002E6161742E612E65455443646C2E2E6E61730000000F41",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"BFA5B112B2B0074360036242BD6203A5004405020000000000405A1A00405A1A",
INIT_01 => X"4300A34300A303004300A3006002100300000007524000000007836000000000",
INIT_02 => X"020300024300A3020040424000A54300A34300A303004300A300800224A50020",
INIT_03 => X"7005B0022311B1BD0440644400620300004402BDE0B0B1B2BF4300A3024300A3",
INIT_04 => X"4202434512B202BDBDE0B0B1BF8400A54005022000000010008443A5BF300262",
INIT_05 => X"024464024003008300620240620213A5000544024060233111B080B1B3B4BF62",
INIT_06 => X"02A500BF050410B0BD004042004202BDE0B0B1B2B3B4BF534343205100426200",
INIT_07 => X"000000E0BD0004B0BF000004A500050405000004A50005040500000400004504",
INIT_08 => X"A560C6A4A3C38404A505C606A560A4A08404A505A560A4A08404A505BD1D9C1C",
INIT_09 => X"AEADACABAAA9A8A7A6A5A4A3A2A1BD0000000000A560C6A4A3C38404A505C606",
INIT_0A => X"BABFB9B8AFAEADACABAAA9A8A7A6A5A4A3A2A10000BB00BB00BA5A1ABFB9B8AF",
INIT_0B => X"00828242038200E0004042008200E000404200820084E0029B401BBD60BB60BB",
INIT_0C => X"402000A540400540400400BFB080B1BD00E08243038200E08242008200E08243",
INIT_0D => X"A542000205402000A542000205402000A502000202420205402000A542000205",
INIT_0E => X"402000A5020002420205402000A5020002420205402000A50200020205402000",
INIT_0F => X"B0B3B4B5B611B1BD000000000000BFBD000000BDE0B0B100BF00000002000202",
INIT_10 => X"B5B6BF3114100400007240004000220040004053424016A2141615000031B2BF",
INIT_11 => X"B120B0BF100400C6201004002044A006B0BF624211B1B102BDBDE0B0B1B2B3B4",
INIT_12 => X"A400650062424302828402008082E043436283430462630343420302BD0004C6",
INIT_13 => X"038000E0606085A400656400E00000636600C3C486006464C5A54462C0A6A4C0",
INIT_14 => X"E4006467600045460062468287E6E2000042E600878246470000C2E047678662",
INIT_15 => X"A20283A2E0A30382000000E00000C6C04060404087E400444764848700470047",
INIT_16 => X"85A2A6C682824302A2830200E085A2A6C682824302A2830200E085A2058283A3",
INIT_17 => X"8243038200E085A500E08582A200E0850000E085A2A6C682824302A2830200E0",
INIT_18 => X"00E0824200820000000000000000E08500E08243420003A08200E085A205A582",
INIT_19 => X"BF93B3BD000000E0824300828242038200E0824300828242038200E082430382",
INIT_1A => X"020202420262020000000202020242026202404040524040A0000480B060B1B2",
INIT_1B => X"0302400400004000203102030300000000024004000040006023021200001202",
INIT_1C => X"05400000A50505400000A50540004240A000BFB0B1BDBDE0B0B1B2B300BF0203",
INIT_1D => X"82C20060C2438683A5400082BDE000B0B1BFBD00B120B0BF05000005400000A5",
INIT_1E => X"BDE000BF000000E0400022E2080020A5A0000500BFA080BD00E000820202E0C5",
INIT_1F => X"0000400082824540008202C000E000820200E0A282A20060A243858300400082",
INIT_20 => X"4000828243A300830040008200C245008200400082824500820040008202C200",
INIT_21 => X"02004022000291BD000000B000B1BF8062B1BFB00243BD8200E08545A3008300",
INIT_22 => X"00BD00B000BF0000040000040000040062024300028000BFB0BD000031004425",
INIT_23 => X"BDE000BF4400426663466400808645658082428000BFBD44E042000060004380",
INIT_24 => X"40004300A382A00060A302C302A3816000074000E700A3C30749200900436404",
INIT_25 => X"B002BF8000B0BFBD0000000000E0648063A4A5808000E042E002434263A50084",
INIT_26 => X"BFB0BDBDE0B0B10011BF8000B1B0B1BFBDBDE0B0B111BF8000A0B0B1BFBDBDE0",
INIT_27 => X"200014103320000052004000021312A080B4BFB0B1B2B3BDBDE042B0BF028000",
INIT_28 => X"840005048400050484000504B000B1BF8400BD0400BDE0B0B1B2B3B4BF000034",
INIT_29 => X"000400620004038400A50405220004118400A510040504008400050484000504",
INIT_2A => X"0004050004A5000405050004050004A5000405050004050004A5000405040004",
INIT_2B => X"BDE000B0B1BF8400A50405A500054402A5000524040004000505000405000405",
INIT_2C => X"656F65003A300A416C0A00616965000061657720694645524E45520D494F5343",
INIT_2D => X"0000000000000000000000000000706500726500656F6500656F6500656F6500",
INIT_2E => X"6469747278004154006462676F62742E0701670000405A1A00405A1A00000000",
INIT_2F => X"00405A1A00405A1A0000000000000000000000000000007362746E4B53627400",
INIT_30 => X"0000007362746E4B536274006469747278004154006462676F62742E07016700",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"0000000E0000000000001700FF17001603170000000000000000040000000400",
INIT_01 => X"0000000000000000000000000016000020049000000000008800000000008020",
INIT_02 => X"1600001600000016000000200400000000000000000000000000001600000420",
INIT_03 => X"00000000170000FF000017000017000004170000000000000000000016000000",
INIT_04 => X"17001601000020FF000000000017041604002017000000000417041600172018",
INIT_05 => X"0016FF0000100016000000A000009E00039E1700800018170000000000000020",
INIT_06 => X"0016030000170000FF000000000040000000000000000000160000880016FF00",
INIT_07 => X"0000000000034000000004171703001700033017170300170003301700031617",
INIT_08 => X"00FF0018000017001600160000FF18001700170000FF18001700170019001700",
INIT_09 => X"0000000000000000000000000000FF010001000200FF00180000170017001600",
INIT_0A => X"00000000000000000000000000000000000000000100D800D800FF7000000000",
INIT_0B => X"00000000FF00000000FF000000000000FF000000006000606000000000000000",
INIT_0C => X"002004160000008000000200008800FF00000010FF0000000000000000000010",
INIT_0D => X"1603FF20000020041603FF200000200416000000000320000020041603002000",
INIT_0E => X"0020041600FF000120000020041600FF000420000020041600FF002000002004",
INIT_0F => X"00000000000000FF000000FF000500FF00000000000000100080200200FF0040",
INIT_10 => X"00000000FF0020022898F8000000000000000010900090000000209880170000",
INIT_11 => X"002800003420020028342002280080000000101718000000FF00000000000000",
INIT_12 => X"30000000001717002000FF1000170000000017000018FF001019FF0000022000",
INIT_13 => X"0000000000000000000000100000FF00000000000000000000FF300000002800",
INIT_14 => X"3800000000000000181700FFFF000000FF000000FFFF0000000040280017FF17",
INIT_15 => X"28000010002800000000000000FF001018100000000000000000002000000000",
INIT_16 => X"0028280000001010100000000000282800000010101000000000002828000018",
INIT_17 => X"0010FF0000000000000000000000000000000000282800000010101000000000",
INIT_18 => X"00000000000000010001000100000000000000100000FF000000000028280000",
INIT_19 => X"000000FF00000000001000000000FF000000001000000000FF0000000010FF00",
INIT_1A => X"0000000120000090000000000000004000000000000080008804009000000000",
INIT_1B => X"0000FF0004000000000000000080002004000000040000000000000010000000",
INIT_1C => X"000020041600000020041600000000888001000000FF00000000000010000000",
INIT_1D => X"0000100018100000000000000000100000000003002000000000000000200416",
INIT_1E => X"0000000010000010FF0000380003200000000038004048FF0000100000000000",
INIT_1F => X"0000000000001000000000000000100000000000000010001810000000000000",
INIT_20 => X"0000000010180000000000000000280000000000000010000000000000000000",
INIT_21 => X"0000FF10000000000328300020000080000000000000FF000000002828000000",
INIT_22 => X"00000400200000040000040000040000000000000080040000FF00FF00040000",
INIT_23 => X"0000000000FFFFFF00000000002030201810FF280400FF100000FF0000000010",
INIT_24 => X"00000000000020040018000000180030FFFF001000384000000000003010101F",
INIT_25 => X"00000080010000FF000200020000FFFF00FF001810100000001010000000FF00",
INIT_26 => X"0000FF00000000100000800100000000FF000000000000800188000000FF0000",
INIT_27 => X"2001FF0000200100000000000000008088000000000000FF0000000000008001",
INIT_28 => X"010200000302000000020000000200000228FF0000000000000000000000FF00",
INIT_29 => X"0340031701400016031600001701010016031620000000010002000001020000",
INIT_2A => X"0203000203A10203000002030002035E02030000020300020312020300400140",
INIT_2B => X"0000100000001704160000160400160016030017020102030000030200020200",
INIT_2C => X"72757600303A00496F48007973760000727600006D4644432044430A4F4C2043",
INIT_2D => X"0000161700001717000016170000697600637600727576007275760072757600",
INIT_2E => X"616E616F742E424F562D756E7400727304006E00000004000000040000001717",
INIT_2F => X"000004000000040000000000000000000000000000000000757475005473612E",
INIT_30 => X"00000000757475005473612E616E616F742E424F562D756E7400727304006E00",
INIT_31 => X"0000000000000000000017000000000000000000000000000000000000000000",
INIT_32 => X"0000171600000000000000001716000000000000000016160000000000000015",
INIT_33 => X"0000000000000000000000000002171700000000000000001717000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"24101C1020180D1A023C4801D8480000C8440000000000000008C40000080000",
INIT_01 => X"06001007001130060700100006F4000A2580120D1A020000100D1A0200001012",
INIT_02 => X"F43008F4010010F400080A25801003001004001130060400100006F40A108025",
INIT_03 => X"01001401500018E000164C01004C00002844002808181C2024000010F4010011",
INIT_04 => X"1000F008001800D8200814181C30AB200800005007000908AB3008141C500004",
INIT_05 => X"20F0FF000D2B00F0000B7F25040803FFB4004400251E2B30001023141C20242B",
INIT_06 => X"002CC81400400010E800260100040028081014181C202400F001032B00F0FF08",
INIT_07 => X"00000008182600101400284010C8004020F4254030C8004010F4254000C8F440",
INIT_08 => X"04FB042A00001000F000D00004FD2A001000100004FD2A00E0001000E0001000",
INIT_09 => X"44403C3834302C2824201C181410983000F0004404FB042A000010001000F000",
INIT_0A => X"5854504C4844403C3834302C2824201C18141000F860125C1058FC0054504C48",
INIT_0B => X"00000001FE00000800FC020004000800FC01000400000800000801681360115C",
INIT_0C => X"04259A74040000254F08531C142518E000080024FD0000080002000000080024",
INIT_0D => X"B430ED000004259AA420F5000004259A940439010010000007259A8400080000",
INIT_0E => X"04259A4805D20000000006259A3804DC0000000006259AC003E600000005259A",
INIT_0F => X"101C2024280014D0000000FF000C14E800000020081418251C25257E07CA0000",
INIT_10 => X"24282C04EC0100BD25250900060000000A000C2424120408200100252560182C",
INIT_11 => X"1825141C4200D501250200C825002501141C2160801F1800E030081014181C20",
INIT_12 => X"2B000800170000002403FC2528000804000400080023F47F24E3FC0020E20001",
INIT_13 => X"0035000800040004000004250800E900000604000400000808F4210C1104230F",
INIT_14 => X"2100080C13001A00250000F8F4040400F3000009F8F4040400072B250D00F400",
INIT_15 => X"04011024080401000000000800E600252525000400040004000810210008000E",
INIT_16 => X"1425040114142427041401000818250401181824270418010008102427101025",
INIT_17 => X"0024C70000080002000800000100080C0000081C2504011C1C2427041C010008",
INIT_18 => X"000800080000008A0084007A0000080C000800240402FB030000080025C00700",
INIT_19 => X"240420D800000008002400000020DF000008002400000010EF0000080024F700",
INIT_1A => X"010C0408000905250A1418401008080009071C080400252825B42025142E181C",
INIT_1B => X"4008F140B40008000A020C1440251025B6040540B4000C000E01010125030114",
INIT_1C => X"0008259A4400030F259A34001A00042525901C1418E0280814181C2025241018",
INIT_1D => X"100125092B211018FF0C000820082514181C203C1825141C0200080104259ACC",
INIT_1E => X"1808001425000225F5001C2101B425FF0B000025142525E80008251C02010800",
INIT_1F => X"26002600041021020008010C0008251C020008000C0125042B210C14000C0004",
INIT_20 => X"060004102121001800060008001321140C001800041021001000050008021000",
INIT_21 => X"0000F32B00100820F425251425181C2509181C140704E00000080C2121001400",
INIT_22 => X"0018B610251400B60000B60800B60400070704000025281410E800F501CF0000",
INIT_23 => X"1808001401F5FFFF01000000082A23232521FF256014E8230801FB0003000025",
INIT_24 => X"0900050000002569002100022D210525F5FF0312301021010D1A020A252326C3",
INIT_25 => X"10081425731014E8007E00530008FFFC01FF01252525080108232BFFFF01F801",
INIT_26 => X"1410E82008141825081C256CFF14181CE020081418081C256C2514181CE01808",
INIT_27 => X"256CFF0108256C0004000D00000D0A252520241014181CD81808FF1014082573",
INIT_28 => X"C427070044270600442702001427181C6025E0000028081014181C202400F108",
INIT_29 => X"30001A40840000488A44000044840000388A34000000016830271F00B4270800",
INIT_2A => X"F82008F32020F020070CF81008F31010F0105F0CF80008F300D0F00013006C00",
INIT_2B => X"20082514181C10AB70000068AB00F40058C80044008400100101070004FC000C",
INIT_2C => X"306E2F003030004E20650030702F0000742F000065002020002020004E415645",
INIT_2D => X"00006810000000000000681000006F2F00302F00336E2F00326E2F00316E2F00",
INIT_2E => X"7469006400744C5245696975652E7468010075000008C4000008000000000000",
INIT_2F => X"0008C40000080000A00002070B000000000000000000000074722E2E41730064",
INIT_30 => X"0000000074722E2E417300647469006400744C5245696975652E746801007500",
INIT_31 => X"D03007012A0001000020900000011E0004000024A00002070B00000000000000",
INIT_32 => X"002070F0030142000100002070D003083801040000D0A00032013000100000D0",
INIT_33 => X"000000000000000053000100000090E003084D00100000D09010030848001000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic